module struct1;
  struct {
    int  a;
    byte b;
  } s1;

  typedef struct {
    int x, y;
  } t_pair;
endmodule // struct1

