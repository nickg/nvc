-- -*- coding: iso-8859-1 -*-
package strings is
    constant s1 : string := "�ngstr�m";
end package;
