architecture a of one is
begin

end architecture;
