architecture a of e is
begin
    f(1, 2, 3 + 5);
    assert x'attr;
end architecture;
