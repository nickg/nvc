module parse1;
  wire [8:0] x, y;
  assign y = x; // + 1;
endmodule // parse1
