-- LCS-2016-082: Empty record
package pack is

    type rec is record
    end record ;

end package ;
