package p is

    type a is (x, y, z);
    type b is ('x', 'y', Z);
    type c is (FOO);
    
end package;
