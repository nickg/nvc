package func is

    function add(x, y : integer; y : in integer) return integer;

    impure function naughty return integer;
    
end package;
