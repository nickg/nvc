package error2 is
    subtype char128 is character range (NUL to DEL);  -- Error
end package;
