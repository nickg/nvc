entity one is
end entity;

entity two is
end two;

entity three is
end entity three;
