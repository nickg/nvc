package pack is
    procedure foo is new bar.all;
end package;
