module union1;
  union { int x; logic y; } u1;
  typedef union { int a; logic b; } t_u2;
endmodule // union1
