PACKAGE p IS

  CONSTANT a : INTEGER := 2#1101#;
  CONSTANT b : INTEGER := 3#20#;
  CONSTANT c : INTEGER := 8#7#;
  CONSTANT d : INTEGER := 10#1234#;
  CONSTANT e : INTEGER := 16#beef01#;
  CONSTANT f : INTEGER := 2#1_0#;
  CONSTANT g : INTEGER := 2:1_0:;
  CONSTANT h : INTEGER := 16#abababab#;
  CONSTANT i : INTEGER := 16#1A#;
  CONSTANT j : INTEGER := 2#1111_1111#;
  CONSTANT k : INTEGER := 16#FF#;
  CONSTANT l : INTEGER := 016#0FF#;
  CONSTANT m : INTEGER := 16#E#E1;
  CONSTANT n : INTEGER := 2#1110_0000#;
  CONSTANT o : REAL    := 16#F.FF#E+2;
  CONSTANT p : REAL    := 2#1.1111_1111_111#E11;
  CONSTANT n : INTEGER := 2:1110_0000:;
  CONSTANT o : REAL    := 16:F.FF:E+2;

END PACKAGE;
