entity issue1060 is
end entity;

architecture test of issue1060 is
begin
end architecture;
