entity bug is
end entity;

architecture a of bug is
begin
  main : process is
  begin
  end;
end;                                    -- Used to hang here
