architecture a of one is
begin

end architecture;

architecture b of one is
begin

end b;

architecture c of one is
begin

end;
