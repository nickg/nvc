entity sub is
    port (
        x : in integer );
end entity;

entity top is
end entity;

architecture test of top is
begin

end architecture;
