architecture a of e is
    signal pos : integer := 64;
    signal neg : integer := -265;
    constant c : integer := 523;
    constant a : string := "hel""lo";
    constant b : string := """quote""";
begin

end architecture;
