architecture a of e is
begin

    x <= a or b;

    x <= 1 when foo
         else 2 when bar
         else 3;
    
end architecture;
