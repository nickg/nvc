-------------------------------------------------------------------------------
--  Copyright (C) 2025  Nick Gasson
--
--  Licensed under the Apache License, Version 2.0 (the "License");
--  you may not use this file except in compliance with the License.
--  You may obtain a copy of the License at
--
--     http://www.apache.org/licenses/LICENSE-2.0
--
--  Unless required by applicable law or agreed to in writing, software
--  distributed under the License is distributed on an "AS IS" BASIS,
--  WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
--  See the License for the specific language governing permissions and
--  limitations under the License.
-------------------------------------------------------------------------------

package body random is

    impure function get_random return t_uint32 is
    begin
        assert false severity failure;
    end function;

    impure function get_random return boolean is
    begin
        return (get_random mod 2) = 0;
    end function;

end package body;
