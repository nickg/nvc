entity ent is
end entity;

architecture a of ent is
begin
  main : process
  begin
    report """""";
    wait;
  end process;
end architecture;
