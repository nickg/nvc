architecture a of e is
begin

    x <= a or b;
    
end architecture;
