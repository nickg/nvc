entity vhpi17 is
end entity;

architecture test of vhpi17 is
begin
end architecture;
