entity assert3 is
begin
    assert (false)
        report "should assert"
        severity note;
end entity assert3;
