hello
`bad
