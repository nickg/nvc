package length is
    -- Seems to be a bug in VHDL-2019 standard
    constant c1 : integer := integer'length;
end package;
