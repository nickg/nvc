-------------------------------------------------------------------------------
--  Copyright (C) 2022  Nick Gasson
--
--  Licensed under the Apache License, Version 2.0 (the "License");
--  you may not use this file except in compliance with the License.
--  You may obtain a copy of the License at
--
--     http://www.apache.org/licenses/LICENSE-2.0
--
--  Unless required by applicable law or agreed to in writing, software
--  distributed under the License is distributed on an "AS IS" BASIS,
--  WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
--  See the License for the specific language governing permissions and
--  limitations under the License.
-------------------------------------------------------------------------------

-------------------------------------------------------------------------------
-- IEEE 1076-2008 section 16.9
-------------------------------------------------------------------------------

context IEEE_BIT_CONTEXT is
    library IEEE;
    use IEEE.NUMERIC_BIT.all;
end context IEEE_BIT_CONTEXT;
