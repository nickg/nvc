package concat is
    constant c1 : bit_vector := "1" & "00";
    constant c2 : string := "xy" & "z";
    constant c3 : bit_vector := '1' & '0';
    constant c4 : string := "fo" & 'o';
end package;
