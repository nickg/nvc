-- -*- coding: iso-8859-1 -*-
entity ����� is
end entity;

architecture ���������� of ����� is
    signal �x�� : bit;
    constant �������������������������������� : integer := 1;
    -- ��������������������������������
    constant ������������������������������ : integer := 2;
begin
end architecture;
