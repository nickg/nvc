package test2 is
  shared variable shared_var : work.test3.t_prot;
end package;
