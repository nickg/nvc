`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XYZ"
`protect encrypt_agent_info = "Foo"
`protect key_keyowner = "Baz", key_keyname = "1235", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
WDaeD6HpPZKvUqmB7Ivy5Ui/FIAwhGoUAogcYLjKWUxEgtiwqmc06LXjNvNbalAzzd6yhHCMgMKx
LspGhgv6XmdjksdgskdlDFDf1qmveCmJc9KH1Yqlhpd1R01IubLx7XzlN9rDwa44wsCcJhayPUDF
bahyL2ThjpwZy6KSCXo=

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 215)
`protect data_block
ZUl11eGlSaTtRJ0hALHF4ND/DxZWOYhtW4EaQDBVpW9aKIUm5tC5AYZFS3JKYbCd3TXgjk6XQ7WX
8gge7eK7U+hWn8pff+iRTPK+L7RstXcOTdVh66EPwVWdjmyPp59duDopJwnJIWH1gJ+0E/0W66KU
m6UCs8b2tN34WadF6E6aP3n1EnfOWf5HyWL/UzUstSa7a9/KrZFanOpl2/pYeEiLpzau7U6ZcJ9/
8zwHfv/PoUCEQiD+/kavwT8L/dZvxNIqTgFzuDUvDkDfA8geLGLV9qvrYJuduajL4Hglz3uQQxAo
D4SpMmUtLi0ru/Sjze7tYn39pEr5quQ4NyGklZAYjlVCp17hLXUY5wA/wmEQzJHTn0Bus8HkMS46
`protect end_protected
