package test_pkg is
  alias alias_t is type_t;
  alias alias_t is type_t;
  constant c : alias_t;
end package;
