-- Missing "library ieee;"
use ieee.math_real.all ;

package RandomPkg is

end RandomPkg ;

package body RandomPkg is
-- Was crash here
end RandomPkg ;
