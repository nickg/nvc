module mod1(one, two, three);
  input one;
  input two;
  output three;
endmodule // mixed1
