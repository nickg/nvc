architecture a of e is
    alias foo is bar;
    alias blah : integer is boo;
begin

end architecture;
