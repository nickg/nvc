module extend(i, o);
  parameter WIDTH;
  input i;
  output [WIDTH-1:0] o;

  assign o = {WIDTH{i}};
endmodule
