package issueH is
    constant c : bit_vector;            -- Should be extern
end package issueH;

package body issueH is
    constant c : bit_vector := "101";
end package body issueH;
