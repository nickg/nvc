entity vhpi5 is
end entity;

architecture test of vhpi5 is
    type rec is record
        x, y : integer;
    end record;

    signal s1 : rec;
begin
end architecture;
