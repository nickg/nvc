architecture a of b is
    type my_int1 is range 0 to 10;
    signal x : my_int1 := 2;
begin

    foo: process is
    begin
    end process;
    
end architecture;
