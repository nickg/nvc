package dummy_pkg;
  wire a;
endpackage : different_name
