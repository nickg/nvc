`resetall                 // OK

module foo;
endmodule // foo
