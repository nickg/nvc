architecture a of e is
begin

    process is
    begin
        x := not y;
        x := abs y;
        x := y ** z;
        x := f(4).z;
    end process;

end architecture;
