architecture a of e is
begin

    x <= guarded y;

    with b select z <= guarded q when others;

end architecture;
