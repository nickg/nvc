architecture a of e is
    alias foo is bar;
    alias blah : integer is boo;

    alias funci is func [integer, boolean return boolean];
    alias proci is proc [integer];
    alias proce is proc [];
    alias funce is func [return integer];
begin

end architecture;
