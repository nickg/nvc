entity e is
end entity;

architecture a of e is
    constant x : integer := 5;

    function f_pure(n : in integer) return integer is
    begin
        return n + 1;
    end function;


begin

    process is
        variable v : integer;
    begin
        v := x;                         -- OK
        x := v;                         -- Error
    end process;

    process is
        constant c : integer;           -- Error
    begin
    end process;

    process is
        constant c : integer := f_pure(5);  -- OK
    begin
    end process;

end architecture;
