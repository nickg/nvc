architecture a of e is
    signal pos : integer := 64;
    signal neg : integer := -265;
    constant c : integer := 523;
    constant a : string := "hel""lo";
    constant b : string := """quote""";
    constant d : integer := 1E3;        -- Integer not real
    constant e : real := 1.234;
    constant f : real := 0.21712;
    constant g : real := 1.4e6;
    constant h : real := 235.1e-2;
begin

end architecture;
