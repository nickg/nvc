entity mre_conversion is
end entity mre_conversion;

architecture arch of mre_conversion is
begin

  mre_conversion_inst: entity work.mre_conversion;

end architecture arch;
