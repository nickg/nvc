entity one is
end entity;

entity two is
end two;

entity three;
end entity three;
