entity noconst is
end noconst;

architecture arch of noconst is
  type map_type is array(bit) of character;
  constant smap : map_type := "";       -- Error
begin
end;
