module lower1;
  wire x, y, z;
  assign z = x & y;
endmodule // lower1
