-- -*- coding: iso-8859-1 -*-
entity ����� is
end entity;

architecture ���������� of ����� is
    signal �x�� : bit;
    constant �������������������������������� : integer := 1;
    -- ��������������������������������
    constant ������������������������������ : integer := 2;

    constant times� :  integer := 3;    -- Error
begin
end architecture;
