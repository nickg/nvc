entity describe1 is
end entity;

architecture test of describe1 is
    signal x : integer := 5;
begin

    b1: block is
        signal y : bit;
    begin
    end block;

end architecture;
