module enum1;
  enum { a, b } [3:0] x;   // OK
  typedef enum { c, d } y;   // OK
endmodule // enum1
