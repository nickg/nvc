package func is

    function add(x, y : integer; y : in integer) return integer;

    impure function naughty return integer;

    function "+"(x, y : integer) return integer;
    
end package;
