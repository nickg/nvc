architecture a of e is
    attribute foo : integer;
    attribute foo of x : signal is 5;
begin
    
end architecture;
