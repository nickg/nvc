module mod1(one, two, three);
  input one;
  input two;
  output three;
  parameter g1;
endmodule // mixed1
