library ieee;
use ieee.std_logic_1164.all;
library work;
entity LogTable_0_10_74_F400_uid60 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(9 downto 0);
          Y : out  std_logic_vector(73 downto 0)   );
end entity;

architecture arch of LogTable_0_10_74_F400_uid60 is
signal TableOut, TableOut_d1 :  std_logic_vector(73 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            TableOut_d1 <=  TableOut;
         end if;
      end process;
  with X select TableOut <=
   "11111111111111101111111111111100000000000000000000000000000000000000000000" when "0000000000",
   "11111111111111101111111111111100000000000000000000000000000000000000000000" when "0000000001",
   "00000000001111110000011111111101010101011001010101100010001001001100110101" when "0000000010",
   "00000000011111110010000000000110101011101010110001000100111011110011100001" when "0000000011",
   "00000000101111110100100000100000000101000100110000101110000000110100101101" when "0000000100",
   "00000000111111111000000001010001100101011000100010110011010101111110010110" when "0000000101",
   "00000001001111111100100010100011010001111000011110001110000111000111011111" when "0000000110",
   "00000001100000000010000100011101010001011000011010110101010000001110000011" when "0000000111",
   "00000001110000001000100111000111101100001110001001111111101010101110110111" when "0000001000",
   "00000010000000010000001010101010101100010001101111001110001001010001100110" when "0000001001",
   "00000010010000011000101111001110011100111101111000111101000100100011100011" when "0000001010",
   "00000010100000100010010100111011001011010000011001011101111100011101010110" when "0000001011",
   "00000010110000101100111011111001000101101010011111111000110000010001010100" when "0000001100",
   "00000011000000111000100100010000011100010001010001010101010001000001001011" when "0000001101",
   "00000011010001000101001110001001100000101110000010001100010000111011001010" when "0000001110",
   "00000011100001010010111001101100100110001110101111100000110011000000001100" when "0000001111",
   "00000011110001100001100111000010000001100110011000100001011101110101110001" when "0000010000",
   "00000100000001110001010110010010001001001101011000010001110100100111110010" when "0000010001",
   "00000100010010000010000111100101010101000001111111011011111001011111111011" when "0000010010",
   "00000100100010010011111011000011111110101000101110001001111100011001010001" when "0000010011",
   "00000100110010100110110000110110100001001100101110001000011001011000100110" when "0000010100",
   "00000101000010111010101001000101011001100000001100110000001001110011001001" when "0000010101",
   "00000101010011001111100011111001000101111100110101011001001011001110100110" when "0000010110",
   "00000101100011100101100001011010000110100100001011110101011111100111000101" when "0000010111",
   "00000101110011111100100001110000111101000000000110110100101001101001000100" when "0000011000",
   "00000110000100010100100101000110001100100011001010101111101000101110011011" when "0000011001",
   "00000110010100101101101011100010011010001001000100011101010111101111100110" when "0000011010",
   "00000110100101000111110101001110001100010111000100001111110001111011000010" when "0000011011",
   "00000110110101100011000010010010001011011100011000111001100001000110111001" when "0000011100",
   "00000111000101111111010010110111000001010010101010111100011000110001111111" when "0000011101",
   "00000111010110011100100111000101011001011110011000000000100001001010111101" when "0000011110",
   "00000111100110111010111111000110000001001111001110010100010101110101101101" when "0000011111",
   "00000111110111011010011011000001100111100000101000010101011011001001001110" when "0000100000",
   "00000111110111011010011011000001100111100000101000010101011011001001001110" when "0000100001",
   "00001000000111111010111011000000111100111010001000100010001110000000101110" when "0000100010",
   "00001000011000011100011111001100110011101111110101010100110001011101010100" when "0000100011",
   "00001000101000111111000111101110000000000010110101000110011101010110010111" when "0000100100",
   "00001000111001100010110100101101010111100001101010011100110001111000110110" when "0000100101",
   "00001001001010000111100110010011110001101000110000011111010011010111000000" when "0000100110",
   "00001001011010101101011100101010000111100010110111010110110001101011101010" when "0000100111",
   "00001001101011010100010111111001010100001001100000110101011111010101111100" when "0000101000",
   "00001001111011111100011000001010010100000101011101001000111011010011111110" when "0000101001",
   "00001010001100100101011101100110000101101111000111110100110001100100010100" when "0000101010",
   "00001010011101001111101000010101101001001111000100110111010101111000010010" when "0000101011",
   "00001010101101111010111000100010000000011110011101110111011100100010000001" when "0000101100",
   "00001010111110100111001110010100001111000111011111011011110100101100000000" when "0000101101",
   "00001011001111010100101001110101011010100101110110101100001000001000001010" when "0000101110",
   "00001011001111010100101001110101011010100101110110101100001000001000001010" when "0000101111",
   "00001011100000000011001011001110101010000111001110111011100100000111011100" when "0000110000",
   "00001011110000110010110010101001000110101011101111011101001111001011111000" when "0000110001",
   "00001100000001100011100000001101111011000110011001100010001111101001000011" when "0000110010",
   "00001100010010010101010100000110010011111101100110100001100110101000110000" when "0000110011",
   "00001100100011001000001110011011011111101011100110001010000011101011000001" when "0000110100",
   "00001100110011111100001111010110101110011110111100111101110100011011000101" when "0000110101",
   "00001101000100110001010111000001010010011011000010111000010100110011111110" when "0000110110",
   "00001101010101100111100101100100011111011000100001111110000011010001101010" when "0000110111",
   "00001101100110011110111011001001101011000101110101010110011101001101011011" when "0000111000",
   "00001101100110011110111011001001101011000101110101010110011101001101011011" when "0000111001",
   "00001101110111010111010111111010001101000111101000010000000111100101110100" when "0000111010",
   "00001110001000010000111011111111011110111001010101001111000111110100100110" when "0000111011",
   "00001110011001001011100111100010111011101101100101100101110000110110111000" when "0000111100",
   "00001110101010000111011010101110000000101110110000110111101000101101010111" when "0000111101",
   "00001110111011000100010101101010001100111111011100100111001010011100110110" when "0000111110",
   "00001111001100000010011000100001000001011010111100001101101000111000101110" when "0000111111",
   "00001111011101000001100011011100000000110101110000111101110110000011011000" when "0001000000",
   "00001111101110000001110110100100101111111110001010010001010011110010001011" when "0001000001",
   "00001111111111000011010010000100110101011100100110000000010001100100110000" when "0001000010",
   "00001111111111000011010010000100110101011100100110000000010001100100110000" when "0001000011",
   "00010000010000000101110110000101111001110100010001000100011100000001011101" when "0001000100",
   "00010000100001001001100010110001100111100011101000000110100010001010010000" when "0001000101",
   "00010000110010001110011000010001101011000100111000010110110101000000010011" when "0001000110",
   "00010001000011010100010110101111110010101110100000110000100101101101011111" when "0001000111",
   "00010001010100011011011110010101101110110011110011001000100110101101111100" when "0001001000",
   "00010001100101100011101111001101010001100101010101100110110100010101010100" when "0001001001",
   "00010001110110101101001001100000001111010001100100001011001001001101100110" when "0001001010",
   "00010001110110101101001001100000001111010001100100001011001001001101100110" when "0001001011",
   "00010010000111110111101101011000011110000101010010011101100011001111110000" when "0001001100",
   "00010010011001000011011010111111110110001100001101101001011101011000000101" when "0001001101",
   "00010010101010010000010010100000010001110001011110100100100010111010100011" when "0001001110",
   "00010010111011011110010100000011101101000000001100000001000000111101101111" when "0001001111",
   "00010011001100101101011111110100000110000011111101001011011010100100101011" when "0001010000",
   "00010011011101111101110101111011011101001001011100010100000100010010100100" when "0001010001",
   "00010011011101111101110101111011011101001001011100010100000100010010100100" when "0001010010",
   "00010011101111001111010110100011110100011110111001100100001011110101001100" when "0001010011",
   "00010100000000100010000001110111010000010100101101111110110000100101010101" when "0001010100",
   "00010100010001110101110111111111110110111101111110101101010001101110100011" when "0001010101",
   "00010100100011001010111001000111110000110001000000011000010110110010000010" when "0001010110",
   "00010100110100100001000101011001001000000111111010101100010111011010011111" when "0001010111",
   "00010101000101111000011100111110001001100001001100001010000111011001011001" when "0001011000",
   "00010101000101111000011100111110001001100001001100001010000111011001011001" when "0001011001",
   "00010101010111010001000000000001000011100000001110000011101011101000000110" when "0001011010",
   "00010101101000101010101110101100000110101101111000100101011101001001111010" when "0001011011",
   "00010101111010000101101001001001100101111001000111001011011111001110000111" when "0001011100",
   "00010110001011100001101111100011110101110111011101000011001101010100000010" when "0001011101",
   "00010110011100111111000010000101001101100101101001111001100110010100110010" when "0001011110",
   "00010110011100111111000010000101001101100101101001111001100110010100110010" when "0001011111",
   "00010110101110011101100000111000000110001000001110110101111001111001100000" when "0001100000",
   "00010110111111111101001100000110111010101100000011100000111101000110110101" when "0001100001",
   "00010111010001011110000011111100001000100110111011011001001011101001001000" when "0001100010",
   "00010111100011000000001000100010001111011000001011010011011010101111001010" when "0001100011",
   "00010111110100100011011010000011110000101001001111001000100011000011111010" when "0001100100",
   "00010111110100100011011010000011110000101001001111001000100011000011111010" when "0001100101",
   "00011000000110000111111000101011010000001110001111110000000110111001111101" when "0001100110",
   "00011000010111101101100100100011010100000110101001000111111001111110011010" when "0001100111",
   "00011000101001010100011101110110100100011101110000101000110000001010111110" when "0001101000",
   "00011000111010111100100100101111101011101011011011101000011000110010000011" when "0001101001",
   "00011001001100100101111001011001010110010100100110001000101011100001110110" when "0001101010",
   "00011001001100100101111001011001010110010100100110001000101011100001110110" when "0001101011",
   "00011001011110010000011011111110010011001011111001110100001100111110100011" when "0001101100",
   "00011001101111111100001100101001010011010010010101001000001111110110000110" when "0001101101",
   "00011010000001101001001011100101001001110111110010101100011000110010011011" when "0001101110",
   "00011010010011010111011000111100101100011011110000110111101010010010100011" when "0001101111",
   "00011010010011010111011000111100101100011011110000110111101010010010100011" when "0001110000",
   "00011010100101000110110100111010110010101101111001100011011110010100110000" when "0001110001",
   "00011010110110110111011111101010010110101110101010001100010011011111011001" when "0001110010",
   "00011011001000101001011001010110010100101111111100000000010011011000100011" when "0001110011",
   "00011011011010011100100010001001101011010101101100011011110111111111010100" when "0001110100",
   "00011011101100010000111010001111011011010110100101110100010101111100101011" when "0001110101",
   "00011011101100010000111010001111011011010110100101110100010101111100101011" when "0001110110",
   "00011011111110000110100001110010100111111100101000010000110001100100011011" when "0001110111",
   "00011100001111111101011000111110010110100101110010110001000100100001110100" when "0001111000",
   "00011100100001110101011111111101101111000100101100100011011010001110001101" when "0001111001",
   "00011100110011101110110110111011111011100001001110101000001000110011000000" when "0001111010",
   "00011100110011101110110110111011111011100001001110101000001000110011000000" when "0001111011",
   "00011101000101101001011110000100001000011001001101100100001100111011011000" when "0001111100",
   "00011101010111100101010101100001100100100001000011100010001110011100110000" when "0001111101",
   "00011101101001100010011101011111100001000100011010100010010100000000100000" when "0001111110",
   "00011101101001100010011101011111100001000100011010100010010100000000100000" when "0001111111",
   "00011101111011100000110110001001010001100110110110111000101011111011111011" when "0010000000",
   "00011110001101100000011111101010001100000100100001111011010000100111001101" when "0010000001",
   "00011110011111100001011010001101101000110010110100111110001110100110010001" when "0010000010",
   "00011110110001100011100101111111000010100001000100011111110010111010100000" when "0010000011",
   "00011110110001100011100101111111000010100001000100011111110010111010100000" when "0010000100",
   "00011111000011100111000011001001110110011001001011100011000111110110110001" when "0010000101",
   "00011111010101101011110001111001100100000000010111011010100110110010011111" when "0010000110",
   "00011111100111110001110010011001101101010111110011100001100101011100000011" when "0010000111",
   "00011111111001111001000100110101110110111101010101100101100101001101100001" when "0010001000",
   "00011111111001111001000100110101110110111101010101100101100101001101100001" when "0010001001",
   "00100000001100000001101001011001100111101100001001111111001011001010001110" when "0010001010",
   "00100000011110001011100000010000101000111101100000011010100111001111000110" when "0010001011",
   "00100000110000010110101001100110100110101001011000110000010001100010100001" when "0010001100",
   "00100000110000010110101001100110100110101001011000110000010001100010100001" when "0010001101",
   "00100001000010100011000101100111001111000111010000001101000100010100100000" when "0010001110",
   "00100001010100110000110100011110010011001110101110101010111001100010100100" when "0010001111",
   "00100001100110111111110110010111100110011000010100011001010010110110101100" when "0010010000",
   "00100001111001010000001011011110111110011110000111110110010010111011111001" when "0010010001",
   "00100001111001010000001011011110111110011110000111110110010010111011111001" when "0010010010",
   "00100010001011100001110100000000010011111100100011110111101111000110011100" when "0010010011",
   "00100010011101110100110000000111100001110011000110000101000000010001001110" when "0010010100",
   "00100010110000001001000000000000100101100100111101100001011010010101010010" when "0010010101",
   "00100010110000001001000000000000100101100100111101100001011010010101010010" when "0010010110",
   "00100011000010011110100011110111011111011001111001100111010001000100010111" when "0010010111",
   "00100011010100110101011011111000010001111110111001010011110001110010001000" when "0010011000",
   "00100011100111001101101000001111000010100110111010100011111000111100011100" when "0010011001",
   "00100011100111001101101000001111000010100110111010100011111000111100011100" when "0010011010",
   "00100011111001100111001001000111111001001011101010000010001011000101100101" when "0010011011",
   "00100100001100000001111110101111000000001110010011000101111000011000000011" when "0010011100",
   "00100100011110011110001001010000100100111000010000000011010010001110010000" when "0010011101",
   "00100100011110011110001001010000100100111000010000000011010010001110010000" when "0010011110",
   "00100100110000111011101000111000110110111011111010101101011010011101000100" when "0010011111",
   "00100101000011011010011101110100001000110101011101001001010011100011010110" when "0010100000",
   "00100101010101111010101000001110101111101011100010110010111001100100101111" when "0010100001",
   "00100101010101111010101000001110101111101011100010110010111001100100101111" when "0010100010",
   "00100101101000011100001000010101000011010000001001110011101011011001100110" when "0010100011",
   "00100101111010111110111110010011011110000001010100101011001100000010000110" when "0010100100",
   "00100110001101100011001010010110011101001001111100001001100011101110001110" when "0010100101",
   "00100110001101100011001010010110011101001001111100001001100011101110001110" when "0010100110",
   "00100110100000001000101100101010100000100010100001011100001000110000100000" when "0010100111",
   "00100110110010101111100101011100001010110010000000101100010111110101000001" when "0010101000",
   "00100111000101010111110100111000000001001110100011110001000011111010101110" when "0010101001",
   "00100111000101010111110100111000000001001110100011110001000011111010101110" when "0010101010",
   "00100111011000000001011011001010101011111110010101010010000101110000110110" when "0010101011",
   "00100111101010101100011000100000110101111000010011111110110010111110000101" when "0010101100",
   "00100111101010101100011000100000110101111000010011111110110010111110000101" when "0010101101",
   "00100111111101011000101101000111001100100101000110010111000100111100000011" when "0010101110",
   "00101000010000000110011001001010100000011111101110100111010111110100111000" when "0010101111",
   "00101000100010110101011100110111100100110110011110110111101001110101100100" when "0010110000",
   "00101000100010110101011100110111100100110110011110110111101001110101100100" when "0010110001",
   "00101000110101100101111000011011001111101011101101101101100011001011111000" when "0010110010",
   "00101001001000010111101100000010011001110110101011000001101111001010101010" when "0010110011",
   "00101001011011001010110111111001111111000100010101001000101110110011110110" when "0010110100",
   "00101001011011001010110111111001111111000100010101001000101110110011110110" when "0010110101",
   "00101001101101111111011100001110111101111000001110001111001101101100000110" when "0010110110",
   "00101010000000110101011001001110010111101101010010001010000001011111111101" when "0010110111",
   "00101010000000110101011001001110010111101101010010001010000001011111111101" when "0010111000",
   "00101010010011101100101111000101010000110110101100011001111101000111001011" when "0010111001",
   "00101010100110100101011110000000110000100000101110100011011111110111001100" when "0010111010",
   "00101010111001011111100110001110000000110001100110111010101001111010011011" when "0010111011",
   "00101010111001011111100110001110000000110001100110111010101001111010011011" when "0010111100",
   "00101011001100011011000111111010001110101010010111100010111110100110100010" when "0010111101",
   "00101011011111011000000011010010101010000111101101100011111101110000010100" when "0010111110",
   "00101011011111011000000011010010101010000111101101100011111101110000010100" when "0010111111",
   "00101011110010010110011000100100100110000010111000110001111101000000110001" when "0011000000",
   "00101100000101010110000111111101011000010010100011101011101010010011011010" when "0011000001",
   "00101100011000010111010001101010011001101011101011101100100000101010110001" when "0011000010",
   "00101100011000010111010001101010011001101011101011101100100000101010110001" when "0011000011",
   "00101100101011011001110101111001000110000010011001110011111000101100101100" when "0011000100",
   "00101100111110011101110100110110111100001010111011100001011101111100111110" when "0011000101",
   "00101100111110011101110100110110111100001010111011100001011101111100111110" when "0011000110",
   "00101101010001100011001110110001011101111010011100000110110010110001100110" when "0011000111",
   "00101101100100101010000011110110010000000111111110001110001100000001010000" when "0011001000",
   "00101101110111110010010100010010111010101101010101110111001110010000110101" when "0011001001",
   "00101101110111110010010100010010111010101101010101110111001110010000110101" when "0011001010",
   "00101110001010111100000000010101001000101000000010101000110110001010110000" when "0011001011",
   "00101110011110000111001000001010100111111010001010011001010101101111001100" when "0011001100",
   "00101110011110000111001000001010100111111010001010011001010101101111001100" when "0011001101",
   "00101110110001010011101100000001001001101011010100001100010000010001110000" when "0011001110",
   "00101111000100100001101100000110100010001001100011100110011110111110010000" when "0011001111",
   "00101111000100100001101100000110100010001001100011100110011110111110010000" when "0011010000",
   "00101111010111110001001000101000101000101010010100011000101000000011010100" when "0011010001",
   "00101111101011000010000001110101010111101011010110011111110010100111010000" when "0011010010",
   "00101111101011000010000001110101010111101011010110011111110010100111010000" when "0011010011",
   "00101111111110010100010111111010101100110011101010011101000001010000001100" when "0011010100",
   "00110000010001101000001011000110101000110100011110000011011101101110011010" when "0011010101",
   "00110000100100111101011011100111001111101010001001011101011111111101010100" when "0011010110",
   "00110000100100111101011011100111001111101010001001011101011111111101010100" when "0011010111",
   "00110000111000010100001001101010101000011101001100101000111010110100001100" when "0011011000",
   "00110001001011101100010101011110111101100011001101001010011001000110010000" when "0011011001",
   "00110001001011101100010101011110111101100011001101001010011001000110010000" when "0011011010",
   "00110001011111000101111111010010011100011111110100011000010101010110101010" when "0011011011",
   "00110001110010100001000111010011010110000101101101111101010111001010101101" when "0011011100",
   "00110001110010100001000111010011010110000101101101111101010111001010101101" when "0011011101",
   "00110010000101111101101101101111111110010111100110110010100000101010001001" when "0011011110",
   "00110010011001011011110010110110101100101001001100010001010111000011101011" when "0011011111",
   "00110010011001011011110010110110101100101001001100010001010111000011101011" when "0011100000",
   "00110010101100111011010110110101111011100000001011111110010001010000101100" when "0011100001",
   "00110011000000011100011001111100001000110101010011101010110111011001111010" when "0011100010",
   "00110011000000011100011001111100001000110101010011101010110111011001111010" when "0011100011",
   "00110011010011111110111100010111110101110101010001110000111110100011111100" when "0011100100",
   "00110011100111100010111110010111100111000001110110000110001011110001000011" when "0011100101",
   "00110011100111100010111110010111100111000001110110000110001011110001000011" when "0011100110",
   "00110011111011001000100000001010000100010010110011001000001001101011010001" when "0011100111",
   "00110100001110101111100001111101111000110110111111100001111100001111111111" when "0011101000",
   "00110100001110101111100001111101111000110110111111100001111100001111111111" when "0011101001",
   "00110100100010011000000100000001110011010101011000001010011101111100100000" when "0011101010",
   "00110100110110000010000110100100100101101110000010011100010010000000111111" when "0011101011",
   "00110100110110000010000110100100100101101110000010011100010010000000111111" when "0011101100",
   "00110101001001101101101001110101000101011011001111000110110111100101011111" when "0011101101",
   "00110101011101011010101110000010001011010010011101011001101001010011010100" when "0011101110",
   "00110101011101011010101110000010001011010010011101011001101001010011010100" when "0011101111",
   "00110101110001001001010011011010110011100101011110101000110101011010111001" when "0011110000",
   "00110110000100111001011010001101111110000011011010001100011010010101001000" when "0011110001",
   "00110110000100111001011010001101111110000011011010001100011010010101001000" when "0011110010",
   "00110110011000101011000010101010101101111001110001111001010011100101011001" when "0011110011",
   "00110110101100011110001101000000001001110101100110110101000011101000001111" when "0011110100",
   "00110110101100011110001101000000001001110101100110110101000011101000001111" when "0011110101",
   "00110111000000010010111001011101011100000100011110100100000110100000111100" when "0011110110",
   "00110111000000010010111001011101011100000100011110100100000110100000111100" when "0011110111",
   "00110111010100001001001000010001110010010101101000110010111001111111010001" when "0011111000",
   "00110111101000000000111001101100011101111011000101011010000111011101001101" when "0011111001",
   "00110111101000000000111001101100011101111011000101011010000111011101001101" when "0011111010",
   "00110111111011111010001101111100110011101010101010111101111100011011010000" when "0011111011",
   "00111000001111110101000101010010001011111111001101101000111110001000110101" when "0011111100",
   "00111000001111110101000101010010001011111111001101101000111110001000110101" when "0011111101",
   "00111000100011110001011111111100000010111001100110100010100101001101011000" when "0011111110",
   "00111000110111101111011110001001111000000001111011100001001110001101001110" when "0011111111",
   "00111000110111101111011110001001111000000001111011100001001110001101001110" when "0100000000",
   "00111001001011101111000000001011001110101000100111011000101100001101010010" when "0100000001",
   "00111001011111110000000110001111101101100111100010100100101010011110100011" when "0100000010",
   "00111001011111110000000110001111101101100111100010100100101010011110100011" when "0100000011",
   "00111001110011110010110000100110111111100011001100001111101010100010111100" when "0100000100",
   "00111001110011110010110000100110111111100011001100001111101010100010111100" when "0100000101",
   "00111010000111110110111111100000110010101011110011110110101100000011000101" when "0100000110",
   "00111010011011111100110011001100111000111110100011001001101011110100110010" when "0100000111",
   "00111010011011111100110011001100111000111110100011001001101011110100110010" when "0100001000",
   "00111010110000000100001011111011001000000110101000101001000111111001000001" when "0100001001",
   "00111011000100001101001001111011011001011110100010100000110101111111110111" when "0100001010",
   "00111011000100001101001001111011011001011110100010100000110101111111110111" when "0100001011",
   "00111011011000010111101101011101101010010001001010000000011010101000010010" when "0100001100",
   "00111011101100100011110110110001111011011010111111010001001110011001011001" when "0100001101",
   "00111011101100100011110110110001111011011010111111010001001110011001011001" when "0100001110",
   "00111100000000110001100110001000010001101011010101101010011111111010100100" when "0100001111",
   "00111100000000110001100110001000010001101011010101101010011111111010100100" when "0100010000",
   "00111100010101000000111011110000110101100101100000100011100000010111011110" when "0100010001",
   "00111100101001010001110111111011110011100010000000100100001001000100111011" when "0100010010",
   "00111100101001010001110111111011110011100010000000100100001001000100111011" when "0100010011",
   "00111100111101100100011010111001011011101111110001010100001000100011101110" when "0100010100",
   "00111101010001111000100100111010000010010101010111101001000101100110001110" when "0100010101",
   "00111101010001111000100100111010000010010101010111101001000101100110001110" when "0100010110",
   "00111101100110001110010110001101111111010010010000010011100111000101110000" when "0100010111",
   "00111101100110001110010110001101111111010010010000010011100111000101110000" when "0100011000",
   "00111101111010100101101111000101101110011111111111001011101111011101010101" when "0100011001",
   "00111110001110111110101111110001101111110011011110111100111010100110110100" when "0100011010",
   "00111110001110111110101111110001101111110011011110111100111010100110110100" when "0100011011",
   "00111110100011011001011000100010100110111110010001010001101101100000111000" when "0100011100",
   "00111110100011011001011000100010100110111110010001010001101101100000111000" when "0100011101",
   "00111110110111110101101001101000111011101111101111011111100110101011101010" when "0100011110",
   "00111111001100010011100011010101011001110110011011110010111110110011001010" when "0100011111",
   "00111111001100010011100011010101011001110110011011110010111110110011001010" when "0100100000",
   "00111111100000110011000101111000110001000001010010111011101001000110111100" when "0100100001",
   "00111111100000110011000101111000110001000001010010111011101001000110111100" when "0100100010",
   "00111111110101010100010001100011110101000000111110011010000011000110111100" when "0100100011",
   "01000000001001110111000110100111011101101001000111001101100011010110100010" when "0100100100",
   "01000000001001110111000110100111011101101001000111001101100011010110100010" when "0100100101",
   "01000000011110011011100101010100100110110001101001000011110111001111101100" when "0100100110",
   "01000000110011000001101101111100010000011000000110001001111111111000101010" when "0100100111",
   "01000000110011000001101101111100010000011000000110001001111111111000101010" when "0100101000",
   "01000001000111101001100000101111011110100000111011011110111110001000011010" when "0100101001",
   "01000001000111101001100000101111011110100000111011011110111110001000011010" when "0100101010",
   "01000001011100010010111101111111011001011000110101101000011110001110001111" when "0100101011",
   "01000001110000111110000101111101001101010110000110001001110011011011000110" when "0100101100",
   "01000001110000111110000101111101001101010110000110001001110011011011000110" when "0100101101",
   "01000010000101101010111000111010001010111001111001011101010100010011111101" when "0100101110",
   "01000010000101101010111000111010001010111001111001011101010100010011111101" when "0100101111",
   "01000010011010011001010111000111100110110001101101010000101000011110000110" when "0100110000",
   "01000010101111001001100000110110111001111000100111100011111000011111101010" when "0100110001",
   "01000010101111001001100000110110111001111000100111100011111000011111101010" when "0100110010",
   "01000011000011111011010110011001100001011000101110001100010001011000101100" when "0100110011",
   "01000011000011111011010110011001100001011000101110001100010001011000101100" when "0100110100",
   "01000011011000101110111000000000111110101100011110111010001100100010001000" when "0100110101",
   "01000011011000101110111000000000111110101100011110111010001100100010001000" when "0100110110",
   "01000011101101100100000101111110110111100000001000000011001101101010010111" when "0100110111",
   "01000100000010011011000000100100110101110011000001110000001000010001000000" when "0100111000",
   "01000100000010011011000000100100110101110011000001110000001000010001000000" when "0100111001",
   "01000100010111010011101000000100100111111001000111101111011110001100111000" when "0100111010",
   "01000100010111010011101000000100100111111001000111101111011110001100111000" when "0100111011",
   "01000100101100001101111100110000000000011100010011101100101001010010001010" when "0100111100",
   "01000101000001001001111110111000110110011101111000001100000001111000001001" when "0100111101",
   "01000101000001001001111110111000110110011101111000001100000001111000001001" when "0100111110",
   "01000101010110000111101110110001000101010111111100001100010100101001000000" when "0100111111",
   "01000101010110000111101110110001000101010111111100001100010100101001000000" when "0101000000",
   "01000101101011000111001100101010101100111110110111001101011001101111110000" when "0101000001",
   "01000101101011000111001100101010101100111110110111001101011001101111110000" when "0101000010",
   "01000110000000001000011000110111110001100010101101111101000000000011011110" when "0101000011",
   "01000110010101001011010011101010011011110000101111101001011110111001110110" when "0101000100",
   "01000110010101001011010011101010011011110000101111101001011110111001110110" when "0101000101",
   "01000110101010001111111101010100111000110100110011111011000001010100101100" when "0101000110",
   "01000110101010001111111101010100111000110100110011111011000001010100101100" when "0101000111",
   "01000110111111010110010110001001011010011010111001010011011101101010100010" when "0101001000",
   "01000110111111010110010110001001011010011010111001010011011101101010100010" when "0101001001",
   "01000111010100011110011110011010010110110000100100010101001100110011111000" when "0101001010",
   "01000111101001101000010110011010001000100110011111010001010100010010110001" when "0101001011",
   "01000111101001101000010110011010001000100110011111010001010100010010110001" when "0101001100",
   "01000111111110110011111110011011001111010001111010011101010110110101000101" when "0101001101",
   "01000111111110110011111110011011001111010001111010011101010110110101000101" when "0101001110",
   "01001000010100000001010110110000001110101110001101010000111110111101011101" when "0101001111",
   "01001000010100000001010110110000001110101110001101010000111110111101011101" when "0101010000",
   "01001000101001010000011111101011101111011110010111101011110111101001111110" when "0101010001",
   "01001000111110100001011001100000011110101110100100100100000110111011011110" when "0101010010",
   "01001000111110100001011001100000011110101110100100100100000110111011011110" when "0101010011",
   "01001001010011110100000100100001001110010101101100011101011110101100000100" when "0101010100",
   "01001001010011110100000100100001001110010101101100011101011110101100000100" when "0101010101",
   "01001001101001001000100001000000110100110110111001001001111000001110111110" when "0101010110",
   "01001001101001001000100001000000110100110110111001001001111000001110111110" when "0101010111",
   "01001001111110011110101111010010001101100011001001110011001110111111111110" when "0101011000",
   "01001010010011110110101111101000011000011010110111101111001111010100100011" when "0101011001",
   "01001010010011110110101111101000011000011010110111101111001111010100100011" when "0101011010",
   "01001010101001010000100010010110011010001111011011111101001110001101010101" when "0101011011",
   "01001010101001010000100010010110011010001111011011111101001110001101010101" when "0101011100",
   "01001010111110101100000111101111011100100100110101001110011111010010010100" when "0101011101",
   "01001010111110101100000111101111011100100100110101001110011111010010010100" when "0101011110",
   "01001011010100001001100000000110101101110011001110111001011110010001000110" when "0101011111",
   "01001011010100001001100000000110101101110011001110111001011110010001000110" when "0101100000",
   "01001011101001101000101011101111100001001000101000011000000001100000100101" when "0101100001",
   "01001011111111001001101010111101001110101010011101010001001011011010110000" when "0101100010",
   "01001011111111001001101010111101001110101010011101010001001011011010110000" when "0101100011",
   "01001100010100101100011110000011010011010111001110001110110000101001011010" when "0101100100",
   "01001100010100101100011110000011010011010111001110001110110000101001011010" when "0101100101",
   "01001100101010010001000101010101010001001000001010011111001001010000001010" when "0101100110",
   "01001100101010010001000101010101010001001000001010011111001001010000001010" when "0101100111",
   "01001100111111110111100001000110101110110010111010000011100011001010101010" when "0101101000",
   "01001100111111110111100001000110101110110010111010000011100011001010101010" when "0101101001",
   "01001101010101011111110001101011011000001011001000101011001100100011101101" when "0101101010",
   "01001101010101011111110001101011011000001011001000101011001100100011101101" when "0101101011",
   "01001101101011001001110111010110111110000100010001011011101100110110110001" when "0101101100",
   "01001110000000110101110010011101010110010011001011000111000011011011011000" when "0101101101",
   "01001110000000110101110010011101010110010011001011000111000011011011011000" when "0101101110",
   "01001110010110100011100011010010011011101111110101001111100011000111010101" when "0101101111",
   "01001110010110100011100011010010011011101111110101001111100011000111010101" when "0101110000",
   "01001110101100010011001010001010001110010111000101111010000010000010001000" when "0101110001",
   "01001110101100010011001010001010001110010111000101111010000010000010001000" when "0101110010",
   "01001111000010000100100111011000110011001100011000001110110101010010110110" when "0101110011",
   "01001111000010000100100111011000110011001100011000001110110101010010110110" when "0101110100",
   "01001111010111110111111011010010010100011011011011101001110000011110101011" when "0101110101",
   "01001111010111110111111011010010010100011011011011101001110000011110101011" when "0101110110",
   "01001111101101101101000110001011000001011010000011111001100000111101011010" when "0101110111",
   "01010000000011100100001000010111001110101001111001101110111101010111010001" when "0101111000",
   "01010000000011100100001000010111001110101001111001101110111101010111010001" when "0101111001",
   "01010000011001011101000010001011010101111010001100011100100001101101110110" when "0101111010",
   "01010000011001011101000010001011010101111010001100011100100001101101110110" when "0101111011",
   "01010000101111010111110011111011110110001001100100000110010001000000111110" when "0101111100",
   "01010000101111010111110011111011110110001001100100000110010001000000111110" when "0101111101",
   "01010001000101010100011101111101010011100111110100100010110101001110110110" when "0101111110",
   "01010001000101010100011101111101010011100111110100100010110101001110110110" when "0101111111",
   "01010001011011010011000000100100010111110111110001001101110110111110001100" when "0110000000",
   "01010001011011010011000000100100010111110111110001001101110110111110001100" when "0110000001",
   "01010001110001010011011100000101110001110001000001101100000110001111101101" when "0110000010",
   "01010001110001010011011100000101110001110001000001101100000110001111101101" when "0110000011",
   "01010010000111010101110000110110010101100001110111000001101110000100011010" when "0110000100",
   "01010010000111010101110000110110010101100001110111000001101110000100011010" when "0110000101",
   "01010010011101011001111111001010111100110001000001111011001100110100110110" when "0110000110",
   "01010010011101011001111111001010111100110001000001111011001100110100110110" when "0110000111",
   "01010010110011100000000111011000100110011111101001101001001011100101111111" when "0110001000",
   "01010011001001101000001001110100010111001011000011101111101110110111001010" when "0110001001",
   "01010011001001101000001001110100010111001011000011101111101110110111001010" when "0110001010",
   "01010011011111110010000110110011011000101110101100101001011011010101111000" when "0110001011",
   "01010011011111110010000110110011011000101110101100101001011011010101111000" when "0110001100",
   "01010011110101111101111110101010111010100110000000111110101001110011010011" when "0110001101",
   "01010011110101111101111110101010111010100110000000111110101001110011010011" when "0110001110",
   "01010100001100001011110001110000010001101110010111110001100101001000000110" when "0110001111",
   "01010100001100001011110001110000010001101110010111110001100101001000000110" when "0110010000",
   "01010100100010011011100000011000111000101000111101011111001110000100000011" when "0110010001",
   "01010100100010011011100000011000111000101000111101011111001110000100000011" when "0110010010",
   "01010100111000101101001010111010001111011100101111110110000000010111001000" when "0110010011",
   "01010100111000101101001010111010001111011100101111110110000000010111001000" when "0110010100",
   "01010101001111000000110001101001111011111000011010100010010101010011000000" when "0110010101",
   "01010101001111000000110001101001111011111000011010100010010101010011000000" when "0110010110",
   "01010101100101010110010100111101101001010100010100110001011111110100101100" when "0110010111",
   "01010101100101010110010100111101101001010100010100110001011111110100101100" when "0110011000",
   "01010101111011101101110101001011001000110100011111101011011110110111101110" when "0110011001",
   "01010101111011101101110101001011001000110100011111101011011110110111101110" when "0110011010",
   "01010110010010000111010010101000010001001010100101100100000010100101100010" when "0110011011",
   "01010110010010000111010010101000010001001010100101100100000010100101100010" when "0110011100",
   "01010110101000100010101101101010111110110111111010000011100001100100111110" when "0110011101",
   "01010110101000100010101101101010111110110111111010000011100001100100111110" when "0110011110",
   "01010110111111000000000110101001010100001111011011000111111011100000101001" when "0110011111",
   "01010110111111000000000110101001010100001111011011000111111011100000101001" when "0110100000",
   "01010111010101011111011101111001011001010111110010111110100110101011111100" when "0110100001",
   "01010111010101011111011101111001011001010111110010111110100110101011111100" when "0110100010",
   "01010111101100000000110011110001011100001101011010110111000110100001001000" when "0110100011",
   "01010111101100000000110011110001011100001101011010110111000110100001001000" when "0110100100",
   "01011000000010100100001000100111110000100100011110101111101001000101110111" when "0110100101",
   "01011000000010100100001000100111110000100100011110101111101001000101110111" when "0110100110",
   "01011000011001001001011100110010110000001011000001111011101010010101000000" when "0110100111",
   "01011000011001001001011100110010110000001011000001111011101010010101000000" when "0110101000",
   "01011000101111110000110000101000111010101011000100100100111011100000110010" when "0110101001",
   "01011000101111110000110000101000111010101011000100100100111011100000110010" when "0110101010",
   "01011001000110011010000100100000110101101100101010000111101110010010010111" when "0110101011",
   "01011001000110011010000100100000110101101100101010000111101110010010010111" when "0110101100",
   "01011001011101000101011000110001001100111000000000101010100010011111101010" when "0110101101",
   "01011001011101000101011000110001001100111000000000101010100010011111101010" when "0110101110",
   "01011001110011110010101101110000110001110111101001010001110110100011101010" when "0110101111",
   "01011001110011110010101101110000110001110111101001010001110110100011101010" when "0110110000",
   "01011010001010100010000011110110011100011010100001010000011010011001001110" when "0110110001",
   "01011010001010100010000011110110011100011010100001010000011010011001001110" when "0110110010",
   "01011010100001010011011011011001001010010110001100010100100101001100001010" when "0110110011",
   "01011010100001010011011011011001001010010110001100010100100101001100001010" when "0110110100",
   "01011010111000000110110100101111111111101000111111110011001110101000011010" when "0110110101",
   "01011010111000000110110100101111111111101000111111110011001110101000011010" when "0110110110",
   "01011011001110111100010000010010000110011100001110110000101100100100010010" when "0110110111",
   "01011011001110111100010000010010000110011100001110110000101100100100010010" when "0110111000",
   "01011011100101110011101110010110101111000110010111001000010110010101111100" when "0110111001",
   "01011011100101110011101110010110101111000110010111001000010110010101111100" when "0110111010",
   "01011011111100101101001111010101010000001101001111110011001111011010100000" when "0110111011",
   "01011011111100101101001111010101010000001101001111110011001111011010100000" when "0110111100",
   "01011100010011101000110011100101000110101000010111101110011011001001100010" when "0110111101",
   "01011100010011101000110011100101000110101000010111101110011011001001100010" when "0110111110",
   "01011100101010100110011011011101110101100011000110000001011100000100110010" when "0110111111",
   "01011100101010100110011011011101110101100011000110000001011100000100110010" when "0111000000",
   "01011101000001100110000111010111000110011110111011000101100001001010010100" when "0111000001",
   "01011101000001100110000111010111000110011110111011000101100001001010010100" when "0111000010",
   "01011101011000100111110111101000101001010101110010101110000100000100001010" when "0111000011",
   "01011101011000100111110111101000101001010101110010101110000100000100001010" when "0111000100",
   "01011101101111101011101100101010010100011100010111010010111011100111001010" when "0111000101",
   "01011101101111101011101100101010010100011100010111010010111011100111001010" when "0111000110",
   "01011110000110110001100110110100000100100100010101111101000110001000101000" when "0111000111",
   "01011110000110110001100110110100000100100100010101111101000110001000101000" when "0111001000",
   "01011110000110110001100110110100000100100100010101111101000110001000101000" when "0111001001",
   "01011110011101111001100110011101111100111110110011110110001111101001011110" when "0111001010",
   "01011110011101111001100110011101111100111110110011110110001111101001011110" when "0111001011",
   "01011110110101000011101100000000000111011110100100011011111000001011011000" when "0111001100",
   "01011110110101000011101100000000000111011110100100011011111000001011011000" when "0111001101",
   "01011111001100001111110111110010110100011010100000110110011110111100100000" when "0111001110",
   "01011111001100001111110111110010110100011010100000110110011110111100100000" when "0111001111",
   "01011111100011011110001010001110011010110000000000010101010111011101000110" when "0111010000",
   "01011111100011011110001010001110011010110000000000010101010111011101000110" when "0111010001",
   "01011111111010101110100011101011011000000101010001101111101101111001110000" when "0111010010",
   "01011111111010101110100011101011011000000101010001101111101101111001110000" when "0111010011",
   "01100000010010000001000100100010010000101011110110001011100000101101011010" when "0111010100",
   "01100000010010000001000100100010010000101011110110001011100000101101011010" when "0111010101",
   "01100000101001010101101101001011101111100010111100101010110101010101110100" when "0111010110",
   "01100000101001010101101101001011101111100010111100101010110101010101110100" when "0111010111",
   "01100001000000101100011110000000100110011001111111000000001110111101110111" when "0111011000",
   "01100001000000101100011110000000100110011001111111000000001110111101110111" when "0111011001",
   "01100001011000000101010111011001101101110010111111101010101101111001100110" when "0111011010",
   "01100001011000000101010111011001101101110010111111101010101101111001100110" when "0111011011",
   "01100001011000000101010111011001101101110010111111101010101101111001100110" when "0111011100",
   "01100001101111100000011001110000000101000101001000111001111111001000111100" when "0111011101",
   "01100001101111100000011001110000000101000101001000111001111111001000111100" when "0111011110",
   "01100010000110111101100101011100110010011111001100111011100011101111000001" when "0111011111",
   "01100010000110111101100101011100110010011111001100111011100011101111000001" when "0111100000",
   "01100010011110011100111010111001000011001010000111010001011000000110000100" when "0111100001",
   "01100010011110011100111010111001000011001010000111010001011000000110000100" when "0111100010",
   "01100010110101111110011010011110001011001011011111010010100011110000110100" when "0111100011",
   "01100010110101111110011010011110001011001011011111010010100011110000110100" when "0111100100",
   "01100011001101100010000100100101100101101000001011110110111010100101011010" when "0111100101",
   "01100011001101100010000100100101100101101000001011110110111010100101011010" when "0111100110",
   "01100011100101000111111001101000110100100110111000001101111000100111011001" when "0111100111",
   "01100011100101000111111001101000110100100110111000001101111000100111011001" when "0111101000",
   "01100011100101000111111001101000110100100110111000001101111000100111011001" when "0111101001",
   "01100011111100101111111010000001100001010010101010000001100010100001100010" when "0111101010",
   "01100011111100101111111010000001100001010010101010000001100010100001100010" when "0111101011",
   "01100100010100011010000110001001011011111101101000100110010100101011010001" when "0111101100",
   "01100100010100011010000110001001011011111101101000100110010100101011010001" when "0111101101",
   "01100100101100000110011110011010011100000011100101011000001011100000011101" when "0111101110",
   "01100100101100000110011110011010011100000011100101011000001011100000011101" when "0111101111",
   "01100101000011110101000011001110100000001100100101100101110000001110010010" when "0111110000",
   "01100101000011110101000011001110100000001100100101100101110000001110010010" when "0111110001",
   "01100101011011100101110100111111101110001111101101001010010101010011111010" when "0111110010",
   "01100101011011100101110100111111101110001111101101001010010101010011111010" when "0111110011",
   "01100101011011100101110100111111101110001111101101001010010101010011111010" when "0111110100",
   "01100101110011011000110100001000010011010101101010110111001110110001011011" when "0111110101",
   "01100101110011011000110100001000010011010101101010110111001110110001011011" when "0111110110",
   "01100110001011001110000001000010100011111011100101101101010010011101001100" when "0111110111",
   "01100110001011001110000001000010100011111011100101101101010010011101001100" when "0111111000",
   "01100110100011000101011100001000111011110101101011100111001101010011010101" when "0111111001",
   "01100110100011000101011100001000111011110101101011100111001101010011010101" when "0111111010",
   "01100110111010111111000101110101111110010010000001010101011010110001110000" when "0111111011",
   "01100110111010111111000101110101111110010010000001010101011010110001110000" when "0111111100",
   "01100110111010111111000101110101111110010010000001010101011010110001110000" when "0111111101",
   "01100111010010111010111110100100010101111011010011101100001100001111011110" when "0111111110",
   "01100111010010111010111110100100010101111011010011101100001100001111011110" when "0111111111",
   "10110110001110010111100110110111000000011110101100001011000011100000101000" when "1000000000",
   "10110110011010010111100000110111001100011110011101001011011101111001100100" when "1000000001",
   "10110110100110010111111110111000100000100010011100011000010000111101110111" when "1000000010",
   "10110110110010011001000000111110010101000100000000011101110101111000000100" when "1000000011",
   "10110110111110011010100111001100000010111010111111110000000000001100111000" when "1000000100",
   "10110111001010011100110001100101000011011101110101111000111011010000011000" when "1000000101",
   "10110111001010011100110001100101000011011101110101111000111011010000011000" when "1000000110",
   "10110111010110011111100000001100110000100001101001101001011101101111011000" when "1000000111",
   "10110111100010100010110011000110100100011010010010101010110100000100110110" when "1000001000",
   "10110111101110100110101010010101111001111010011111010001100001110100011000" when "1000001001",
   "10110111111010101011000101111110001100010011111010010001111010100001111010" when "1000001010",
   "10111000000110110000000110000010110111010111010000110101110010011111111000" when "1000001011",
   "10111000010010110101101010100111010111010100011000010011100111101100001010" when "1000001100",
   "10111000011110111011110011101111001000111010010100000111000011010101011001" when "1000001101",
   "10111000011110111011110011101111001000111010010100000111000011010101011001" when "1000001110",
   "10111000101011000010100001011101101001010111011011101010110100100001011101" when "1000001111",
   "10111000110111001001110011110110010110011001100000010100000100001110010111" when "1000010000",
   "10111001000011010001101010111100101110001101110011001111000011000111010010" when "1000010001",
   "10111001001111011010000110110100001111100001001011011101010001100110110111" when "1000010010",
   "10111001011011100011000111100000011001100000001011110101000010100000110010" when "1000010011",
   "10111001100111101100101101000100101011110111001001000010011000101100001100" when "1000010100",
   "10111001110011110110110111100100100110110010001111101001100000001001000011" when "1000010101",
   "10111001110011110110110111100100100110110010001111101001100000001001000011" when "1000010110",
   "10111010000000000001100111000011101010111101101010001010100010111010011101" when "1000010111",
   "10111010001100001100111011100101011001100101100111000110111010010000000001" when "1000011000",
   "10111010011000011000110101001101010100010110011111000111111100011000110100" when "1000011001",
   "10111010100100100101010011111110111101011100111011000111000111011010010100" when "1000011010",
   "10111010110000110010010111111101110111100101111010010111101001100101111000" when "1000011011",
   "10111010111101000000000001001101100101111110111000110001100111100111101001" when "1000011100",
   "10111010111101000000000001001101100101111110111000110001100111100111101001" when "1000011101",
   "10111011001001001110001111110001101100010101110100111110100001001001101000" when "1000011110",
   "10111011010101011101000011101101101110111001010110100111010100000110000101" when "1000011111",
   "10111011100001101100011101000101010010011000110100100011111111000100100000" when "1000100000",
   "10111011101101111100011011111011111100000100011011001100100011011100001010" when "1000100001",
   "10111011111010001101000000010101010001101101010010101011100111011000000110" when "1000100010",
   "10111100000110011110001010010100111001100101100101010010011000010111111100" when "1000100011",
   "10111100000110011110001010010100111001100101100101010010011000010111111100" when "1000100100",
   "10111100010010101111111001111110011010100000100101101110001110101001010000" when "1000100101",
   "10111100011111000010001111010101011011110010110101011111110001110101100010" when "1000100110",
   "10111100101011010101001010011101100101010010001011010011011111100000100111" when "1000100111",
   "10111100110111101000101011011010011111010101111001011011110011110100000000" when "1000101000",
   "10111101000011111100110010001111110010110110110100001100110100110011001110" when "1000101001",
   "10111101010000010001011111000001001001001111011000011001100000110101101110" when "1000101010",
   "10111101010000010001011111000001001001001111011000011001100000110101101110" when "1000101011",
   "10111101011100100110110001110010001100011011110001110010100000100011000000" when "1000101100",
   "10111101101000111100101010100110100110111010000001100110011100101101111110" when "1000101101",
   "10111101110101010011001001100010000011101010000101000011111000101011111101" when "1000101110",
   "10111110000001101010001110101000001110001101111011111100110001100100111101" when "1000101111",
   "10111110001110000001111001111100110010101001101111001011100010111010010000" when "1000110000",
   "10111110001110000001111001111100110010101001101111001011100010111010010000" when "1000110001",
   "10111110011010011010001011100011011101100011110111011001110001000000100110" when "1000110010",
   "10111110100110110011000011011111111100000101000011101000011001101011110100" when "1000110011",
   "10111110110011001100100001110101111011111000011111111001101011101001010001" when "1000110100",
   "10111110111111100110100110101001001011001011111011111100100101000111011000" when "1000110101",
   "10111111001100000001010001111101011000101111110001111001111010000111110110" when "1000110110",
   "10111111001100000001010001111101011000101111110001111001111010000111110110" when "1000110111",
   "10111111011000011100100011110110010011110111001101000011000010111011000110" when "1000111000",
   "10111111100100111000011100010111101100011000010000100010010011000011001101" when "1000111001",
   "10111111110001010100111011100101010010101011111110001100111001011100101011" when "1000111010",
   "10111111111101110010000001100010110111101110011101010110101010001011111101" when "1000111011",
   "10111111111101110010000001100010110111101110011101010110101010001011111101" when "1000111100",
   "11000000001010001111101110010100001100111111000001100111010010001110011010" when "1000111101",
   "11000000010110101110000001111101000100100000010001110001010101101101110011" when "1000111110",
   "11000000100011001100111100100001010000111000001110101010111001010101010110" when "1000111111",
   "11000000101111101100011110000100100101010000011010000111110111000111111011" when "1001000000",
   "11000000111100001100100110101010110101010101111101110101111111010110101001" when "1001000001",
   "11000000111100001100100110101010110101010101111101110101111111010110101001" when "1001000010",
   "11000001001000101101010110010111110101011001110010011010100101110111101011" when "1001000011",
   "11000001010101001110101101001111011010010000100110010001111100011101000001" when "1001000100",
   "11000001100001110000101011010101011001010011000100110000011010101011011001" when "1001000101",
   "11000001101110010011010000101101101000011101111101000101010011110001010000" when "1001000110",
   "11000001101110010011010000101101101000011101111101000101010011110001010000" when "1001000111",
   "11000001111010110110011101011011111110010010001001011111011010111110011100" when "1001001000",
   "11000010000111011010010001100100010001110100110110010011010110111100111001" when "1001001001",
   "11000010010011111110101101001010011010101111101001000011100100101011001000" when "1001001010",
   "11000010100000100011110000010010010001010000100111101010001010011001100010" when "1001001011",
   "11000010101101001001011010111111101110001010011111100100011011001011001110" when "1001001100",
   "11000010101101001001011010111111101110001010011111100100011011001011001110" when "1001001101",
   "11000010111001101111101101010110101010110100101101000000001011011100000010" when "1001001110",
   "11000011000110010110100111011011000001001011100010001010110111001100110010" when "1001001111",
   "11000011010010111110001001010000101011110000001110100010011010010111101000" when "1001010000",
   "11000011011111100110010010111011100101101001000110000111111011101110000010" when "1001010001",
   "11000011011111100110010010111011100101101001000110000111111011101110000010" when "1001010010",
   "11000011101100001111000100011111101010100001101000110100001011000010101100" when "1001010011",
   "11000011111000111000011110000000110110101010101001101101110011000000111111" when "1001010100",
   "11000100000101100010011111100011000110111010010110100001011111010100111101" when "1001010101",
   "11000100010010001101001001001010011000101100011110111011110111100101110001" when "1001010110",
   "11000100010010001101001001001010011000101100011110111011110111100101110001" when "1001010111",
   "11000100011110111000011010111010101010000010011100000101001111100101100111" when "1001011000",
   "11000100101011100100010100110111111001100011010111111111001101011001111101" when "1001011001",
   "11000100111000010000110111000110000110011100010101000100000101111111000100" when "1001011010",
   "11000101000100111110000001101001010000100000010101101000010000101010001011" when "1001011011",
   "11000101000100111110000001101001010000100000010101101000010000101010001011" when "1001011100",
   "11000101010001101011110100100101011000001000100011011101010010001101111000" when "1001011101",
   "11000101011110011010001111111110011110010100010111010111000000000011111110" when "1001011110",
   "11000101101011001001010011111000100100101001100000110010011100000001001010" when "1001011111",
   "11000101101011001001010011111000100100101001100000110010011100000001001010" when "1001100000",
   "11000101110111111001000000010111101101010100001101011110101001010110010000" when "1001100001",
   "11000110000100101001010101011111111011000111010001000111011011100011001100" when "1001100010",
   "11000110010001011010010011010101010001011100001101000001111111100000011010" when "1001100011",
   "11000110011110001011111001111011110100010011010111111011011111100011001011" when "1001100100",
   "11000110011110001011111001111011110100010011010111111011011111100011001011" when "1001100101",
   "11000110101010111110001001010111101000010100000101101001100011000001100011" when "1001100110",
   "11000110110111110001000001101100110010101100101110111100101001111011010001" when "1001100111",
   "11000111000100100100100010111111011001010010111001010100100101001100100110" when "1001101000",
   "11000111010001011000101101010011100010100011011110110110101100010000100110" when "1001101001",
   "11000111010001011000101101010011100010100011011110110110101100010000100110" when "1001101010",
   "11000111011110001101100000101101010101100010110110000110010000011000101101" when "1001101011",
   "11000111101011000010111101010000111001111100111001111110101110011110111110" when "1001101100",
   "11000111110111111001000011000010011000000101010001101111111111111001101000" when "1001101101",
   "11000111110111111001000011000010011000000101010001101111111111111001101000" when "1001101110",
   "11001000000100101111110010000101111000110111011000111100101010110101110000" when "1001101111",
   "11001000010001100111001010011111100101110110100111011010010010111111110111" when "1001110000",
   "11001000011110011111001100010011101001001110011001010011101011000000110010" when "1001110001",
   "11001000011110011111001100010011101001001110011001010011101011000000110010" when "1001110010",
   "11001000101011010111110111100110001101110010010111001101000111010110000100" when "1001110011",
   "11001000111000010001001100011011011110111110011110001010110011001100111000" when "1001110100",
   "11001001000101001011001010110111101000110111000111111001001000000110100011" when "1001110101",
   "11001001010010000101110010111110111000001001010010110111001000101110110000" when "1001110110",
   "11001001010010000101110010111110111000001001010010110111001000101110110000" when "1001110111",
   "11001001011111000001000100110101011010001010101010100010111111101010100110" when "1001111000",
   "11001001101011111101000000011111011100111001101111101000100010101001000010" when "1001111001",
   "11001001111000111001100110000001001110111110000000010001111010111100011100" when "1001111010",
   "11001001111000111001100110000001001110111110000000010001111010111100011100" when "1001111011",
   "11001010000101110110110101011110111111101000000000011010010011100110001101" when "1001111100",
   "11001010010010110100101110111100111110110001100010000010101101111100100000" when "1001111101",
   "11001010011111110011010010011111011100111101101101101000111101010011100110" when "1001111110",
   "11001010011111110011010010011111011100111101101101101000111101010011100110" when "1001111111",
   "11001010101100110010100000001010101011011001001010100000101010010011011010" when "1010000000",
   "11001010111001110010011000000010111011111010000111001110011110100011000100" when "1010000001",
   "11001011000110110010111010001100100001000000100010000101011001010011011110" when "1010000010",
   "11001011000110110010111010001100100001000000100010000101011001010011011110" when "1010000011",
   "11001011010011110100000110101011101101110110010001100110001101110011011000" when "1010000100",
   "11001011100000110101111101100100110110001111001101000001001011110110010011" when "1010000101",
   "11001011101101111000011110111100001110101001010100111001110011011001001000" when "1010000110",
   "11001011101101111000011110111100001110101001010100111001110011011001001000" when "1010000111",
   "11001011111010111011101010110110001100001100111011101100110011101110011010" when "1010001000",
   "11001100000111111111100001010111000100101100101110011000010110111101101000" when "1010001001",
   "11001100010101000100000010100011001110100101111101000110011010011111110001" when "1010001010",
   "11001100010101000100000010100011001110100101111101000110011010011111110001" when "1010001011",
   "11001100100010001001001110011111000001000000100011111001010101000101000100" when "1010001100",
   "11001100101111001111000101001110110011101111010011011010101011001110111000" when "1010001101",
   "11001100111100010101100110110110111111001111111001101100010010101001101100" when "1010001110",
   "11001100111100010101100110110110111111001111111001101100010010101001101100" when "1010001111",
   "11001101001001011100110011011011111100101011001010111011100101010011000110" when "1010010000",
   "11001101010110100100101011000010000101110101001010010111000100110111110110" when "1010010001",
   "11001101100011101101001101101101110101001101010011000110001111010110101001" when "1010010010",
   "11001101100011101101001101101101110101001101010011000110001111010110101001" when "1010010011",
   "11001101110000110110011011100011100101111110100001000011100101010100001000" when "1010010100",
   "11001101111110000000010100100111110011111111011001111001000010101101010000" when "1010010101",
   "11001110001011001010111000111110111011110010010101111110101010110100111011" when "1010010110",
   "11001110001011001010111000111110111011110010010101111110101010110100111011" when "1010010111",
   "11001110011000010110001000101101011010100101101001011011101000001010101001" when "1010011000",
   "11001110100101100010000011110111101110010011101101001001100000110111110000" when "1010011001",
   "11001110110010101110101010100010010101100011000111111010000000100001001011" when "1010011010",
   "11001110110010101110101010100010010101100011000111111010000000100001001011" when "1010011011",
   "11001110111111111011111100110001101111100110110111011110110111111100000000" when "1010011100",
   "11001111001101001001111010101010011100011110011001110100010011110011010011" when "1010011101",
   "11001111011010011000100100010000111100110101110110001101101010101101111101" when "1010011110",
   "11001111011010011000100100010000111100110101110110001101101010101101111101" when "1010011111",
   "11001111100111100111111001101001110010000110000110100100100011100011100100" when "1010100000",
   "11001111110100110111111010111001011110010101000000101010010100101111100100" when "1010100001",
   "11001111110100110111111010111001011110010101000000101010010100101111100100" when "1010100010",
   "11010000000010001000101000000100100100010101011111011011111101010010010010" when "1010100011",
   "11010000001111011010000001001111100111100111101100011000011000001111100010" when "1010100100",
   "11010000011100101100000110011111001100011001001000111001001011011011001100" when "1010100101",
   "11010000011100101100000110011111001100011001001000111001001011011011001100" when "1010100110",
   "11010000101001111110110111110111110111100100110111101101110010000011100101" when "1010100111",
   "11010000110111010010010101011110001110110011100110011001000100001010110010" when "1010101000",
   "11010000110111010010010101011110001110110011100110011001000100001010110010" when "1010101001",
   "11010001000100100110011111010110111000011011110110110001011011011111100110" when "1010101010",
   "11010001010001111011010101100110011011100010001000100011010110100111010001" when "1010101011",
   "11010001011111010000111000010001011111111001000010110110011011001001100100" when "1010101100",
   "11010001011111010000111000010001011111111001000010110110011011001001100100" when "1010101101",
   "11010001101100100111000111011100101110000001011101110100110111110000111010" when "1010101110",
   "11010001111001111110000011001100101111001010101100010101100110110000100101" when "1010101111",
   "11010010000111010101101011100110001101010010100101101000110010000011011011" when "1010110000",
   "11010010000111010101101011100110001101010010100101101000110010000011011011" when "1010110001",
   "11010010010100101110000000101101110011000101101111000110111001010101011100" when "1010110010",
   "11010010100010000111000010101000001011111111100110000010011011001011011100" when "1010110011",
   "11010010100010000111000010101000001011111111100110000010011011001011011100" when "1010110100",
   "11010010101111100000110001011010000100001010101001011100000001111011101110" when "1010110101",
   "11010010111100111011001101001000001000100000100011111001010101001011011000" when "1010110110",
   "11010011001010010110010101110111000110101010010101011110010000100100000001" when "1010110111",
   "11010011001010010110010101110111000110101010010101011110010000100100000001" when "1010111000",
   "11010011010111110010001011101011101101000000011101101001000000110101110110" when "1010111001",
   "11010011100101001110101110101010101010101011000101010000100111111010101001" when "1010111010",
   "11010011100101001110101110101010101010101011000101010000100111111010101001" when "1010111011",
   "11010011110010101011111110111000101111100010001000100110001000101110010000" when "1010111100",
   "11010100000000001001111100011010101100001101100001011000011011110001100001" when "1010111101",
   "11010100000000001001111100011010101100001101100001011000011011110001100001" when "1010111110",
   "11010100001101101000100111010101010010000101010000111010101101001100111100" when "1010111111",
   "11010100011011000111111111101101010011010001101010001101100101001000110011" when "1011000000",
   "11010100101000101000000101100111100010101011011100001010111011010000100000" when "1011000001",
   "11010100101000101000000101100111100010101011011100001010111011010000100000" when "1011000010",
   "11010100110110001000111001001000110011111011111011110100010110010111010010" when "1011000011",
   "11010101000011101010011010010101111011011101001110100100011000110101000110" when "1011000100",
   "11010101000011101010011010010101111011011101001110100100011000110101000110" when "1011000101",
   "11010101010001001100101001010011101110011010010100100010011010110010001010" when "1011000110",
   "11010101011110101111100110000111000010101111010010111001010010111000100101" when "1011000111",
   "11010101011110101111100110000111000010101111010010111001010010111000100101" when "1011001000",
   "11010101101100010011010000110100101111001001011110010000101110100011100000" when "1011001001",
   "11010101111001110111101001100001101011000111100101001001011010100011010111" when "1011001010",
   "11010110000111011100110000010010101110111001111010011011111100101111101100" when "1011001011",
   "11010110000111011100110000010010101110111001111010011011111100101111101100" when "1011001100",
   "11010110010101000010100101001100110011100010011111111010011111111110101001" when "1011001101",
   "11010110100010101001001000010100110010110101010000110101010010111011010000" when "1011001110",
   "11010110100010101001001000010100110010110101010000110101010010111011010000" when "1011001111",
   "11010110110000010000011001101111100111011000001100100001111010110011010000" when "1011010000",
   "11010110111101111000011001100010001100100011100001000101011010110110001110" when "1011010001",
   "11010110111101111000011001100010001100100011100001000101011010110110001110" when "1011010010",
   "11010111001011100001000111110001011110100001110110000001010001011111100011" when "1011010011",
   "11010111011001001010100100100010011010010000010111000011001100000101100001" when "1011010100",
   "11010111011001001010100100100010011010010000010111000011001100000101100001" when "1011010101",
   "11010111100110110100101111111001111101011110111110110111110010000111110010" when "1011010110",
   "11010111110100011111101001111101000110110000100010000000001000111000010000" when "1011010111",
   "11010111110100011111101001111101000110110000100010000000001000111000010000" when "1011011000",
   "11011000000010001011010010110000110101011010111001101010010000011001010011" when "1011011001",
   "11011000001111110111101010011010001001100111001110101100011010101100111010" when "1011011010",
   "11011000011101100100110000111110000100010010000100100011011110010000100101" when "1011011011",
   "11011000011101100100110000111110000100010010000100100011011110010000100101" when "1011011100",
   "11011000101011010010100110100001100111001011100100010100000100100010000011" when "1011011101",
   "11011000111001000001001011001001110100110111100111101110110101101001100010" when "1011011110",
   "11011000111001000001001011001001110100110111100111101110110101101001100010" when "1011011111",
   "11011001000110110000011110111011110000101110000100010111100010000110010011" when "1011100000",
   "11011001010100100000100001111100011110111010110110101111001011011010110010" when "1011100001",
   "11011001010100100000100001111100011110111010110110101111001011011010110010" when "1011100010",
   "11011001100010010001010100010001000100011110001101100001001100110101110100" when "1011100011",
   "11011001110000000010110101111110100111001100110100110011100100110111001011" when "1011100100",
   "11011001110000000010110101111110100111001100110100110011100100110111001011" when "1011100101",
   "11011001111101110101000111001010001101110000000001011010000000101101011101" when "1011100110",
   "11011010001011101000000111111000111111100101111100001100001010101100001010" when "1011100111",
   "11011010001011101000000111111000111111100101111100001100001010101100001010" when "1011101000",
   "11011010011001011011111000010000000101000001101101011110111100011001000111" when "1011101001",
   "11011010100111010000011000010100100111001011101000100000110101110000011101" when "1011101010",
   "11011010100111010000011000010100100111001011101000100000110101110000011101" when "1011101011",
   "11011010110101000101101000001011110000000001010110111001011001111111010001" when "1011101100",
   "11011011000010111011100111111010101010010110000100001011110011010100110100" when "1011101101",
   "11011011000010111011100111111010101010010110000100001011110011010100110100" when "1011101110",
   "11011011010000110010010111100110100001110010101001011100011110101011000100" when "1011101111",
   "11011011011110101001110111010100100010110101111000111010000000000111100100" when "1011110000",
   "11011011011110101001110111010100100010110101111000111010000000000111100100" when "1011110001",
   "11011011101100100010000111001001111010110100101001101001000001010101110000" when "1011110010",
   "11011011111010011011000111001011110111111010000011010011011010111100101110" when "1011110011",
   "11011011111010011011000111001011110111111010000011010011011010111100101110" when "1011110100",
   "11011100001000010100110111011111101001000111101001111010101001110010010000" when "1011110101",
   "11011100010110001111011000001010011110010101101001101101010001001101111101" when "1011110110",
   "11011100010110001111011000001010011110010101101001101101010001001101111101" when "1011110111",
   "11011100100100001010101001010001101000010011000010111111101011011111010000" when "1011111000",
   "11011100110010000110101010111010011000100101110110001000001001001001011000" when "1011111001",
   "11011100110010000110101010111010011000100101110110001000001001001001011000" when "1011111010",
   "11011101000000000011011101001010000001101011001111011110000000101001011111" when "1011111011",
   "11011101001110000001000000000101110110110111110011011100001111001010100000" when "1011111100",
   "11011101001110000001000000000101110110110111110011011100001111001010100000" when "1011111101",
   "11011101011011111111010011110011001100010111101010100111001011101011110000" when "1011111110",
   "11011101101001111110011000010111010111001110101101110101101101011110110001" when "1011111111",
   "11011101101001111110011000010111010111001110101101110101101101011110110001" when "1100000000",
   "11011101110111111110001101110111101101011000110010011101100111000010000110" when "1100000001",
   "11011110000101111110110100011001100101101001110110100011010110011110100010" when "1100000010",
   "11011110000101111110110100011001100101101001110110100011010110011110100010" when "1100000011",
   "11011110010100000000001100000010010111101110001101001101001100101101000100" when "1100000100",
   "11011110010100000000001100000010010111101110001101001101001100101101000100" when "1100000101",
   "11011110100010000010010100110111011100001010101010111001101100001100001101" when "1100000110",
   "11011110110000000101001110111110001100011100110001111001100000101011100011" when "1100000111",
   "11011110110000000101001110111110001100011100110001111001100000101011100011" when "1100001000",
   "11011110111110001000111010011100000010111010111110101100110000110101001110" when "1100001001",
   "11011111001100001101010111010110011010110100110100100011101010111100111010" when "1100001010",
   "11011111001100001101010111010110011010110100110100100011101010111100111010" when "1100001011",
   "11011111011010010010100101110010110000010011001010000010101101111100110100" when "1100001100",
   "11011111101000011000100101110110100000011000010101101010001111101001011101" when "1100001101",
   "11011111101000011000100101110110100000011000010101101010001111101001011101" when "1100001110",
   "11011111110110011111010111100111001001000000011010100001100001100101001000" when "1100001111",
   "11100000000100100110111011001010001001000001010101000101010101011101000111" when "1100010000",
   "11100000000100100110111011001010001001000001010101000101010101011101000111" when "1100010001",
   "11100000010010101111010000100101000000001011000111111010000010011010010001" when "1100010010",
   "11100000010010101111010000100101000000001011000111111010000010011010010001" when "1100010011",
   "11100000100000111000010111111101001111001000001000100001001100001111110100" when "1100010100",
   "11100000101111000010010001011000010111011101001100010010101101110011001100" when "1100010101",
   "11100000101111000010010001011000010111011101001100010010101101110011001100" when "1100010110",
   "11100000111101001100111100111011111011101001110101011001100111101000001101" when "1100010111",
   "11100001001011011000011010101101011111001000011111110100010100001101110101" when "1100011000",
   "11100001001011011000011010101101011111001000011111110100010100001101110101" when "1100011001",
   "11100001011001100100101010110010100110001110101110011000100010110111011001" when "1100011010",
   "11100001100111110001101101010000110110001101010111111010111010011111011101" when "1100011011",
   "11100001100111110001101101010000110110001101010111111010111010011111011101" when "1100011100",
   "11100001110101111111100010001101110101010000110100011010000101100001010110" when "1100011101",
   "11100001110101111111100010001101110101010000110100011010000101100001010110" when "1100011110",
   "11100010000100001110001001101111001010100001001010001101101000000111001010" when "1100011111",
   "11100010010010011101100011111010011110000010011011011000100001111010100101" when "1100100000",
   "11100010010010011101100011111010011110000010011011011000100001111010100101" when "1100100001",
   "11100010100000101101110000110101011000110100110010111111011100100110111010" when "1100100010",
   "11100010101110111110110000100101100100110100110010100010101000011011110010" when "1100100011",
   "11100010101110111110110000100101100100110100110010100010101000011011110010" when "1100100100",
   "11100010111101010000100011010000101100111011011111011011101000000000000000" when "1100100101",
   "11100011001011100011001000111100011100111110110000011110101100100100101100" when "1100100110",
   "11100011001011100011001000111100011100111110110000011110101100100100101100" when "1100100111",
   "11100011011001110110100001101110100001110001011011100000000100001001011110" when "1100101000",
   "11100011011001110110100001101110100001110001011011100000000100001001011110" when "1100101001",
   "11100011101000001010101101101100101001000011100010111100111010100010101000" when "1100101010",
   "11100011110110011111101100111100100001100010100011101000001110110010111100" when "1100101011",
   "11100011110110011111101100111100100001100010100011101000001110110010111100" when "1100101100",
   "11100100000100110101011111100011111010111001100010011011011110001011011100" when "1100101101",
   "11100100010011001100000101101000100101110001011010001011000110000011010101" when "1100101110",
   "11100100010011001100000101101000100101110001011010001011000110000011010101" when "1100101111",
   "11100100100001100011011111010000010011110001001001011110111101111011110001" when "1100110000",
   "11100100100001100011011111010000010011110001001001011110111101111011110001" when "1100110001",
   "11100100101111111011101100100000110111011110000000101110101011000010011100" when "1100110010",
   "11100100111110010100101101100000000100011011110000000001101110100111110100" when "1100110011",
   "11100100111110010100101101100000000100011011110000000001101110100111110100" when "1100110100",
   "11100101001100101110100010010011101111001100110101010011110000011101000001" when "1100110101",
   "11100101001100101110100010010011101111001100110101010011110000011101000001" when "1100110110",
   "11100101011011001001001011000001101101010010101010011100100110101111010001" when "1100110111",
   "11100101101001100100100111101111110101001101110011011100011100110101110010" when "1100111000",
   "11100101101001100100100111101111110101001101110011011100011100110101110010" when "1100111001",
   "11100101111000000000111000100011111110011110001100101011111010001001001000" when "1100111010",
   "11100110000110011101111101100100000001100011011001010000001010011010010110" when "1100111011",
   "11100110000110011101111101100100000001100011011001010000001010011010010110" when "1100111100",
   "11100110010100111011110110110101110111111100110001010011001001000001001101" when "1100111101",
   "11100110010100111011110110110101110111111100110001010011001001000001001101" when "1100111110",
   "11100110100011011010100100011111011100001001110000011111110000011001101100" when "1100111111",
   "11100110110001111010000110100110101001101010000100100010001111001000110010" when "1101000000",
   "11100110110001111010000110100110101001101010000100100010001111001000110010" when "1101000001",
   "11100111000000011010011101010001011100111101111011101100100100000001101111" when "1101000010",
   "11100111000000011010011101010001011100111101111011101100100100000001101111" when "1101000011",
   "11100111001110111011101000100101110011100110010011011111000010100101001101" when "1101000100",
   "11100111011101011101101000101001101100000101000111010101000001010100010100" when "1101000101",
   "11100111011101011101101000101001101100000101000111010101000001010100010100" when "1101000110",
   "11100111101100000000011101100011000101111101011111010101110011010010010010" when "1101000111",
   "11100111101100000000011101100011000101111101011111010101110011010010010010" when "1101001000",
   "11100111111010100100000111011000000001110011111111001001101110001111110001" when "1101001001",
   "11101000001001001000100110001110100001001110110100110011011110111011101110" when "1101001010",
   "11101000001001001000100110001110100001001110110100110011011110111011101110" when "1101001011",
   "11101000010111101101111010001100100110110110000111101101101100110101111010" when "1101001100",
   "11101000010111101101111010001100100110110110000111101101101100110101111010" when "1101001101",
   "11101000100110010100000011011000010110010100000111101100101111000000001110" when "1101001110",
   "11101000110100111011000001110111110100010101011100000100110011001100000000" when "1101001111",
   "11101000110100111011000001110111110100010101011100000100110011001100000000" when "1101010000",
   "11101001000011100010110101110001000110101001010010110100011001000001101110" when "1101010001",
   "11101001000011100010110101110001000110101001010010110100011001000001101110" when "1101010010",
   "11101001010010001011011111001010010100000001101111110011000010100001001110" when "1101010011",
   "11101001100000110100111110001001100100010011111100000100011011011010010011" when "1101010100",
   "11101001100000110100111110001001100100010011111100000100011011011010010011" when "1101010101",
   "11101001101111011111010010110101000000011000010101001111111000111100111101" when "1101010110",
   "11101001101111011111010010110101000000011000010101001111111000111100111101" when "1101010111",
   "11101001111110001010011101010010110010001010111100111100010011100010000100" when "1101011000",
   "11101010001100110110011101101001000100101011101000010000011011101101011010" when "1101011001",
   "11101010001100110110011101101001000100101011101000010000011011101101011010" when "1101011010",
   "11101010011011100011010011111110000011111110001111010111101100001010100100" when "1101011011",
   "11101010011011100011010011111110000011111110001111010111101100001010100100" when "1101011100",
   "11101010101010010001000000010111111101001010111101001011011010000111001110" when "1101011101",
   "11101010111000111111100010111100111110011110011111000000100101101101100010" when "1101011110",
   "11101010111000111111100010111100111110011110011111000000100101101101100010" when "1101011111",
   "11101011000111101110111011110011010111001010010100011010001100000010000011" when "1101100000",
   "11101011000111101110111011110011010111001010010100011010001100000010000011" when "1101100001",
   "11101011010110011111001011000001010111100100111110111111111100001001100001" when "1101100010",
   "11101011010110011111001011000001010111100100111110111111111100001001100001" when "1101100011",
   "11101011100101010000010000101101010001001010010010011001110000111011000011" when "1101100100",
   "11101011110100000010001100111101010110011011100100001111110001000100010110" when "1101100101",
   "11101011110100000010001100111101010110011011100100001111110001000100010110" when "1101100110",
   "11101100000010110100111111110111111010111111111100001110110111000101101010" when "1101100111",
   "11101100000010110100111111110111111010111111111100001110110111000101101010" when "1101101000",
   "11101100010001101000101001100011010011100100100100010010000010101100101001" when "1101101001",
   "11101100100000011101001010000101110101111100111000110000010101010100110111" when "1101101010",
   "11101100100000011101001010000101110101111100111000110000010101010100110111" when "1101101011",
   "11101100101111010010100001100101111001000010111000101111011011010110011010" when "1101101100",
   "11101100101111010010100001100101111001000010111000101111011011010110011010" when "1101101101",
   "11101100111110001000110000001001110100110111010110011011000011101011000100" when "1101101110",
   "11101100111110001000110000001001110100110111010110011011000011101011000100" when "1101101111",
   "11101101001100111111110101111000000010100010000111100001000111010011010110" when "1101110000",
   "11101101011011110111110010110110111100010010010101110010100010100101011000" when "1101110001",
   "11101101011011110111110010110110111100010010010101110010100010100101011000" when "1101110010",
   "11101101101010110000100111001100111101011110101111101001000001110000010010" when "1101110011",
   "11101101101010110000100111001100111101011110101111101001000001110000010010" when "1101110100",
   "11101101111001101010010011000000100010100101111000110001100010011111100100" when "1101110101",
   "11101110001000100100110110011000001001001110011010111011101100001010000110" when "1101110110",
   "11101110001000100100110110011000001001001110011010111011101100001010000110" when "1101110111",
   "11101110010111100000010001011010010000000111010110101110000000011001111010" when "1101111000",
   "11101110010111100000010001011010010000000111010110101110000000011001111010" when "1101111001",
   "11101110100110011100100100001101010111001000010100011111000101111001110110" when "1101111010",
   "11101110100110011100100100001101010111001000010100011111000101111001110110" when "1101111011",
   "11101110110101011001101110110111111111010001110101010011101110110111010100" when "1101111100",
   "11101111000100010111110001100000101010101101100100000001111101000110110101" when "1101111101",
   "11101111000100010111110001100000101010101101100100000001111101000110110101" when "1101111110",
   "11101111010011010110101100001101111100101110100110011001000101011011000010" when "1101111111",
   "11101111010011010110101100001101111100101110100110011001000101011011000010" when "1110000000",
   "11101111100010010110011111000110011001110001101110001110110011111110010011" when "1110000001",
   "11101111100010010110011111000110011001110001101110001110110011111110010011" when "1110000010",
   "11101111110001010111001010010000100111011101101010110001010011011111110011" when "1110000011",
   "11110000000000011000101101110011001100100011011001111110011001000101111011" when "1110000100",
   "11110000000000011000101101110011001100100011011001111110011001000101111011" when "1110000101",
   "11110000001111011011001001110100110000111110011001111111110110011000001110" when "1110000110",
   "11110000001111011011001001110100110000111110011001111111110110011000001110" when "1110000111",
   "11110000011110011110011110011011111101110100111010101100110011110100000110" when "1110001000",
   "11110000011110011110011110011011111101110100111010101100110011110100000110" when "1110001001",
   "11110000101101100010101011101111011101011000001111010000010101000000001111" when "1110001010",
   "11110000101101100010101011101111011101011000001111010000010101000000001111" when "1110001011",
   "11110000111100100111110001110101111011000100111111110101001000110011001001" when "1110001100",
   "11110001001011101101110000110110000011100011011011010110100111000010011100" when "1110001101",
   "11110001001011101101110000110110000011100011011011010110100111000010011100" when "1110001110",
   "11110001011010110100101000110110100100100111101001010110111101110000111000" when "1110001111",
   "11110001011010110100101000110110100100100111101001010110111101110000111000" when "1110010000",
   "11110001101001111100011001111110001101010001111011111010101111110010000001" when "1110010001",
   "11110001101001111100011001111110001101010001111011111010101111110010000001" when "1110010010",
   "11110001111001000101000100010011101101101111000001101001100110011011001010" when "1110010011",
   "11110001111001000101000100010011101101101111000001101001100110011011001010" when "1110010100",
   "11110010001000001110100111111101110111011000010111110100011000011010010001" when "1110010101",
   "11110010010111011001000101000011011100110100011100100000100111101011100110" when "1110010110",
   "11110010010111011001000101000011011100110100011100100000100111101011100110" when "1110010111",
   "11110010100110100100011011101011010001110111000000111001011000001000100000" when "1110011000",
   "11110010100110100100011011101011010001110111000000111001011000001000100000" when "1110011001",
   "11110010110101110000101011111100001011100001011011100101100001001010000001" when "1110011010",
   "11110010110101110000101011111100001011100001011011100101100001001010000001" when "1110011011",
   "11110011000100111101110101111101000000000010111011000011011011111010110010" when "1110011100",
   "11110011000100111101110101111101000000000010111011000011011011111010110010" when "1110011101",
   "11110011010100001011111001110100100110111000111000001010010000010100110000" when "1110011110",
   "11110011100011011010110111101001111000101111001000110000100010100111111110" when "1110011111",
   "11110011100011011010110111101001111000101111001000110000100010100111111110" when "1110100000",
   "11110011110010101010101111100011101111100000010010011000100011101000010011" when "1110100001",
   "11110011110010101010101111100011101111100000010010011000100011101000010011" when "1110100010",
   "11110100000001111011100001101001000110010101111101000010000101100001000111" when "1110100011",
   "11110100000001111011100001101001000110010101111101000010000101100001000111" when "1110100100",
   "11110100010001001101001110000000111001101001000110000001110111001110010110" when "1110100101",
   "11110100010001001101001110000000111001101001000110000001110111001110010110" when "1110100110",
   "11110100100000011111110100110010000111000010010010111110101000011011111001" when "1110100111",
   "11110100101111110011010110000011101101011010000100110011111000001100000110" when "1110101000",
   "11110100101111110011010110000011101101011010000100110011111000001100000110" when "1110101001",
   "11110100111111000111110001111100101100111001001010111010010000001000000110" when "1110101010",
   "11110100111111000111110001111100101100111001001010111010010000001000000110" when "1110101011",
   "11110101001110011101001000100100000110111000110110010101101110011100101011" when "1110101100",
   "11110101001110011101001000100100000110111000110110010101101110011100101011" when "1110101101",
   "11110101011101110011011010000000111110000011001101001001100000100111101011" when "1110101110",
   "11110101011101110011011010000000111110000011001101001001100000100111101011" when "1110101111",
   "11110101101101001010100110011010010110010011011101110001110000111010110101" when "1110110000",
   "11110101101101001010100110011010010110010011011101110001110000111010110101" when "1110110001",
   "11110101111100100010101101110111010100110110010010100011001000111001100001" when "1110110010",
   "11110101111100100010101101110111010100110110010010100011001000111001100001" when "1110110011",
   "11110110001011111011110000011111000000001010000101010000001010110111111101" when "1110110100",
   "11110110011011010101101110011000011111111111010010110100100100100011011111" when "1110110101",
   "11110110011011010101101110011000011111111111010010110100100100100011011111" when "1110110110",
   "11110110101010110000100111101010111101011000101111000110011100111011110101" when "1110110111",
   "11110110101010110000100111101010111101011000101111000110011100111011110101" when "1110111000",
   "11110110111010001100011100011101100010101011111000101101011111100111000010" when "1110111001",
   "11110110111010001100011100011101100010101011111000101101011111100111000010" when "1110111010",
   "11110111001001101001001100110111011011100001001101000000000111101001101100" when "1110111011",
   "11110111001001101001001100110111011011100001001101000000000111101001101100" when "1110111100",
   "11110111011001000110111000111111110100110100011100000110101100001110110111" when "1110111101",
   "11110111011001000110111000111111110100110100011100000110101100001110110111" when "1110111110",
   "11110111101000100101100000111101111100110100111101000100110001001011011110" when "1110111111",
   "11110111101000100101100000111101111100110100111101000100110001001011011110" when "1111000000",
   "11110111111000000101000100111001000011000110000010001000011101101001111100" when "1111000001",
   "11111000000111100101100100111000011000011111001100111111111011001100000111" when "1111000010",
   "11111000000111100101100100111000011000011111001100111111111011001100000111" when "1111000011",
   "11111000010111000111000001000011001111001100100011010100111111010001111100" when "1111000100",
   "11111000010111000111000001000011001111001100100011010100111111010001111100" when "1111000101",
   "11111000100110101001011001100000111010101111000011001111000001110100110101" when "1111000110",
   "11111000100110101001011001100000111010101111000011001111000001110100110101" when "1111000111",
   "11111000110110001100101110011000101111111100110111111011000010101000001011" when "1111001000",
   "11111000110110001100101110011000101111111100110111111011000010101000001011" when "1111001001",
   "11111001000101110000111111110010000101000001101110011010000000010000101100" when "1111001010",
   "11111001000101110000111111110010000101000001101110011010000000010000101100" when "1111001011",
   "11111001010101010110001101110100010001011111001010010101100010100101000111" when "1111001100",
   "11111001010101010110001101110100010001011111001010010101100010100101000111" when "1111001101",
   "11111001100100111100011000100110101110001100111010111010111011001011111110" when "1111001110",
   "11111001100100111100011000100110101110001100111010111010111011001011111110" when "1111001111",
   "11111001110100100011100000010000110101011001001111111100011110001010100110" when "1111010000",
   "11111001110100100011100000010000110101011001001111111100011110001010100110" when "1111010001",
   "11111010000100001011100100111010000010101001001110111001010101011011011000" when "1111010010",
   "11111010000100001011100100111010000010101001001110111001010101011011011000" when "1111010011",
   "11111010010011110100100110101001110010111001001000001011110001000001011000" when "1111010100",
   "11111010100011011110100101100111100100011100101100011101110110110001000011" when "1111010101",
   "11111010100011011110100101100111100100011100101100011101110110110001000011" when "1111010110",
   "11111010110011001001100001111010110110111111100010000100110011100110100010" when "1111010111",
   "11111010110011001001100001111010110110111111100010000100110011100110100010" when "1111011000",
   "11111011000010110101011011101011001011100101011010100010110001000011001011" when "1111011001",
   "11111011000010110101011011101011001011100101011010100010110001000011001011" when "1111011010",
   "11111011010010100010010011000000000100101010101000001111010001001100110000" when "1111011011",
   "11111011010010100010010011000000000100101010101000001111010001001100110000" when "1111011100",
   "11111011100010010000001000000001000110000100010100000110010011101010000100" when "1111011101",
   "11111011100010010000001000000001000110000100010100000110010011101010000100" when "1111011110",
   "11111011110001111110111010110101110101000000110011011110000101111001110000" when "1111011111",
   "11111011110001111110111010110101110101000000110011011110000101111001110000" when "1111100000",
   "11111100000001101110101011100101111000000111111110000011100001100000110001" when "1111100001",
   "11111100000001101110101011100101111000000111111110000011100001100000110001" when "1111100010",
   "11111100010001011111011010011000110111011011100011111101011010101111100010" when "1111100011",
   "11111100010001011111011010011000110111011011100011111101011010101111100010" when "1111100100",
   "11111100100001010001000111010110011100010111100011110110100001111101101000" when "1111100101",
   "11111100100001010001000111010110011100010111100011110110100001111101101000" when "1111100110",
   "11111100110001000011110010100110010001110010100001001110011010011100110110" when "1111100111",
   "11111100110001000011110010100110010001110010100001001110011010011100110110" when "1111101000",
   "11111101000000110111011100010000000011111101111010110001001001000101101101" when "1111101001",
   "11111101000000110111011100010000000011111101111010110001001001000101101101" when "1111101010",
   "11111101010000101100000100011011100000100110100000110101111101100000101010" when "1111101011",
   "11111101010000101100000100011011100000100110100000110101111101100000101010" when "1111101100",
   "11111101100000100001101011010000010110110100101100000100111000001111111110" when "1111101101",
   "11111101100000100001101011010000010110110100101100000100111000001111111110" when "1111101110",
   "11111101110000011000010000110110010111001100110100000011010000011111111111" when "1111101111",
   "11111101110000011000010000110110010111001100110100000011010000011111111111" when "1111110000",
   "11111110000000001111110101010101010011101111100110000111011100000011110010" when "1111110001",
   "11111110000000001111110101010101010011101111100110000111011100000011110010" when "1111110010",
   "11111110010000001000011000110100111111111010011100010011011100000110010110" when "1111110011",
   "11111110010000001000011000110100111111111010011100010011011100000110010110" when "1111110100",
   "11111110100000000001111011011101010000100111110100010110110001011000011111" when "1111110101",
   "11111110100000000001111011011101010000100111110100010110110001011000011111" when "1111110110",
   "11111110101111111100011101010101111100001111100110110111011010100101101100" when "1111110111",
   "11111110101111111100011101010101111100001111100110110111011010100101101100" when "1111111000",
   "11111110111111110111111110100110111010100111011110100001111111011010111111" when "1111111001",
   "11111110111111110111111110100110111010100111011110100001111111011010111111" when "1111111010",
   "11111111001111110100011111011000000101000011001111100001001011001011101100" when "1111111011",
   "11111111001111110100011111011000000101000011001111100001001011001011101100" when "1111111100",
   "11111111011111110001111111110001010110010101001110111100011001100001110110" when "1111111101",
   "11111111011111110001111111110001010110010101001110111100011001100001110110" when "1111111110",
   "11111111101111110000011111111010101010101110101010011101111000001000100000" when "1111111111",
   "--------------------------------------------------------------------------" when others;
    Y <= TableOut_d1;
end architecture;

-------------------------------------------------------------------------------

entity bigcase is
end entity;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

architecture test of bigcase is
    signal clk, rst : std_logic;
    signal X        : std_logic_vector(9 downto 0);
    signal Y        : std_logic_vector(73 downto 0);
begin

    LogTable_0_10_74_F400_uid60_1: entity work.LogTable_0_10_74_F400_uid60
        port map (
            clk => clk,
            rst => rst,
            X   => X,
            Y   => Y );

    p1: process is
        variable ctr : unsigned(9 downto 0);
    begin
        for rep in 1 to 10000 loop
            for i in 1 to 2**9 - 1 loop
                X <= std_logic_vector(ctr);
                ctr := ctr + 1;
                wait for 1 ns;
            end loop;
        end loop;
        wait;
    end process;

end architecture;
