entity vhpi10 is
    generic (
        g0 : integer := 42
        );
end entity;

architecture test of vhpi10 is
begin

end architecture;
