package bitstring is

    constant x : t := X"1234";
    constant y : t := O"1234";
    constant z : t := X"ab";
    constant b : t := B"101";
    
end package;
