library ieee ;

entity issue731 is
end entity ;

architecture arch of issue731 is

    signal bi : ieee.numeric_bit.unsigned(186 downto 0) := d"98234789237429847239487234982347239487239487238947492783" ;

begin

    tb : process
    begin
        assert ieee.numeric_bit.to_string(bi) = "1000000000110011110011110100101110010110101110101110010010011111001001000000111010010001101101101100010111111110011101110101101011111100001110111010010110111101111010100000101001110101111";
        wait;
    end process ;

end architecture ;
