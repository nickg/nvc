entity slow1 is
end entity;

architecture test of slow1 is
    signal finalAdderIn1_bh119 :  bit_vector(60 downto 0);
    signal heap_bh119_w60_3_d1 :  bit;
    signal heap_bh119_w61_2_d1 :  bit;
    signal heap_bh119_w62_1_d1 :  bit;
    signal heap_bh119_w58_3_d1 :  bit;
    signal heap_bh119_w59_2_d1 :  bit;
    signal heap_bh119_w54_4_d2 :  bit;
    signal heap_bh119_w55_3_d2 :  bit;
    signal heap_bh119_w52_4_d2 :  bit;
    signal heap_bh119_w53_3_d2 :  bit;
    signal heap_bh119_w54_3_d2 :  bit;
    signal heap_bh119_w50_4_d2 :  bit;
    signal heap_bh119_w51_3_d2 :  bit;
    signal heap_bh119_w52_3_d2 :  bit;
    signal heap_bh119_w48_4_d2 :  bit;
    signal heap_bh119_w49_3_d2 :  bit;
    signal heap_bh119_w50_3_d2 :  bit;
    signal heap_bh119_w46_4_d2 :  bit;
    signal heap_bh119_w47_3_d2 :  bit;
    signal heap_bh119_w48_3_d2 :  bit;
    signal heap_bh119_w44_4_d2 :  bit;
    signal heap_bh119_w45_3_d2 :  bit;
    signal heap_bh119_w46_3_d2 :  bit;
    signal heap_bh119_w42_4_d2 :  bit;
    signal heap_bh119_w43_3_d2 :  bit;
    signal heap_bh119_w44_3_d2 :  bit;
    signal heap_bh119_w40_4_d2 :  bit;
    signal heap_bh119_w41_3_d2 :  bit;
    signal heap_bh119_w42_3_d2 :  bit;
    signal heap_bh119_w38_4_d2 :  bit;
    signal heap_bh119_w39_3_d2 :  bit;
    signal heap_bh119_w40_3_d2 :  bit;
    signal heap_bh119_w36_4_d2 :  bit;
    signal heap_bh119_w37_3_d2 :  bit;
    signal heap_bh119_w38_3_d2 :  bit;
    signal heap_bh119_w34_4_d2 :  bit;
    signal heap_bh119_w35_3_d2 :  bit;
    signal heap_bh119_w36_3_d2 :  bit;
    signal heap_bh119_w32_4_d2 :  bit;
    signal heap_bh119_w33_3_d2 :  bit;
    signal heap_bh119_w34_3_d2 :  bit;
    signal heap_bh119_w30_4_d2 :  bit;
    signal heap_bh119_w31_3_d2 :  bit;
    signal heap_bh119_w32_3_d2 :  bit;
    signal heap_bh119_w28_4_d2 :  bit;
    signal heap_bh119_w29_3_d2 :  bit;
    signal heap_bh119_w30_3_d2 :  bit;
    signal heap_bh119_w26_4_d2 :  bit;
    signal heap_bh119_w27_3_d2 :  bit;
    signal heap_bh119_w28_3_d2 :  bit;
    signal heap_bh119_w24_4_d2 :  bit;
    signal heap_bh119_w25_3_d2 :  bit;
    signal heap_bh119_w26_3_d2 :  bit;
    signal heap_bh119_w22_4_d2 :  bit;
    signal heap_bh119_w23_3_d2 :  bit;
    signal heap_bh119_w24_3_d2 :  bit;
    signal heap_bh119_w20_4_d2 :  bit;
    signal heap_bh119_w21_3_d2 :  bit;
    signal heap_bh119_w22_3_d2 :  bit;
    signal heap_bh119_w18_4_d2 :  bit;
    signal heap_bh119_w19_3_d2 :  bit;
    signal heap_bh119_w20_3_d2 :  bit;
    signal heap_bh119_w14_4_d2 :  bit;
    signal heap_bh119_w15_3_d2 :  bit;
    signal heap_bh119_w16_3_d2 :  bit;
    signal heap_bh119_w12_3_d2 :  bit;
    signal heap_bh119_w13_3_d2 :  bit;
    signal heap_bh119_w14_3_d2 :  bit;
    signal heap_bh119_w16_4_d2 :  bit;
    signal heap_bh119_w17_3_d2 :  bit;
    signal heap_bh119_w18_3_d2 :  bit;
    signal heap_bh119_w6_0_d2 :  bit;
    signal heap_bh119_w7_0_d2 :  bit;
    signal heap_bh119_w8_0_d2 :  bit;
    signal heap_bh119_w9_0_d2 :  bit;
    signal heap_bh119_w10_0_d2 :  bit;
    signal heap_bh119_w11_0_d2 :  bit;
begin
    -- From flopoco.vhdl
    finalAdderIn1_bh119 <= "0" & '0' & '0' & '0' & heap_bh119_w62_1_d1 & '0' & '0' & '0' & '0' & '0' & '0' & heap_bh119_w55_3_d2 & heap_bh119_w54_3_d2 & heap_bh119_w53_3_d2 & heap_bh119_w52_3_d2 & heap_bh119_w51_3_d2 & heap_bh119_w50_3_d2 & heap_bh119_w49_3_d2 & heap_bh119_w48_3_d2 & heap_bh119_w47_3_d2 & heap_bh119_w46_3_d2 & heap_bh119_w45_3_d2 & heap_bh119_w44_3_d2 & heap_bh119_w43_3_d2 & heap_bh119_w42_3_d2 & heap_bh119_w41_3_d2 & heap_bh119_w40_3_d2 & heap_bh119_w39_3_d2 & heap_bh119_w38_3_d2 & heap_bh119_w37_3_d2 & heap_bh119_w36_3_d2 & heap_bh119_w35_3_d2 & heap_bh119_w34_3_d2 & heap_bh119_w33_3_d2 & heap_bh119_w32_3_d2 & heap_bh119_w31_3_d2 & heap_bh119_w30_3_d2 & heap_bh119_w29_3_d2 & heap_bh119_w28_3_d2 & heap_bh119_w27_3_d2 & heap_bh119_w26_3_d2 & heap_bh119_w25_3_d2 & heap_bh119_w24_3_d2 & heap_bh119_w23_3_d2 & heap_bh119_w22_3_d2 & heap_bh119_w21_3_d2 & heap_bh119_w20_3_d2 & heap_bh119_w19_3_d2 & heap_bh119_w18_3_d2 & heap_bh119_w17_3_d2 & heap_bh119_w16_3_d2 & heap_bh119_w15_3_d2 & heap_bh119_w14_3_d2 & heap_bh119_w13_3_d2 & '0' & heap_bh119_w11_0_d2 & heap_bh119_w10_0_d2 & heap_bh119_w9_0_d2 & heap_bh119_w8_0_d2 & heap_bh119_w7_0_d2 & heap_bh119_w6_0_d2;
end architecture;
