module mod1(i1, o1);
  input [7:0] i1;
  output [3:0] o1;
endmodule // mod1
