package p is

    constant a : integer := 2#1101#;
    constant b : integer := 3#20#;
    constant c : integer := 8#7#;
    constant d : integer := 10#1234#;
    constant e : integer := 16#beef01#;
    constant f : integer := 2#1_0#;
    constant g : integer := 2:1_0:;

end package;
