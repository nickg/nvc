module error1;
  localparam foo bar = 0; // Error
endmodule // error1
