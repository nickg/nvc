architecture a of b is
begin

    -- Wait statements
    process is
    begin
        wait for 1 ns;
    end process;
    
end architecture;
