entity examine1 is
end entity;

library ieee;
use ieee.std_logic_1164.all;

architecture test of examine1 is
    signal x : integer := 5;
    signal y : integer;
    signal a : std_logic := '1';
    signal b : std_logic_vector(3 downto 0) := "01XU";
begin

end architecture;
