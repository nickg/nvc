-- -*- coding: utf-8 -*-
package test is
    constant Åxyzß : bit := '1';          -- Warning
end package;
