entity one is
end entity;

architecture a of one is
    signal x    : integer;
    signal y, z : integer := 7;
begin

end architecture;

architecture b of one is
begin

end b;

architecture c of one is
begin

end;
