package test is
  constant C_ZERO                    : bit_vector(4 downto 0) := 5d"0";
  constant C_ONE                     : bit_vector(4 downto 0) := 5d"1";
  constant C_TWO                     : bit_vector(4 downto 0) := 5d"2";
  constant C_THREE                   : bit_vector(4 downto 0) := 5d"3";
  constant C_TWENTY                  : bit_vector(4 downto 0) := 5d"20";
end package test;
