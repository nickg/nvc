entity one is
end entity;

entity two is
end two;

entity three is
end entity three;

entity four is
    port (
        a : in integer;
        b : out bit;
        c : inout integer;
        d : buffer bit );
end entity;
