context test_context is
end context;

-------------------------------------------------------------------------------

library test_context;
use test_context.test_context.all;      -- Error

entity test is
end entity test;
