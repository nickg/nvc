architecture a of e is
    attribute foo : integer;
begin
    
end architecture;
