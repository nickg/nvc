module Name;
endmodule // Name

module name;
endmodule // name
