`timescale 1ps/1ps
module clkbuf (input i, output o);

  assign o = i;

endmodule // clkmux
