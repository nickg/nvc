architecture a of e is
    signal pos : integer := 64;
    signal neg : integer := -265;
begin

end architecture;
