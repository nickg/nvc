architecture a of e is
    attribute foo : integer;
    attribute foo of x : signal is 5;
    attribute foo of x : component is 5;
begin

end architecture;
