architecture a of b is
    type my_int is range 0 to 100;
    signal x : my_int := 2;
begin

end architecture;
