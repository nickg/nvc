module sub(o);
  parameter i = 0;
  output [7:0] o;
  assign o = i;
endmodule // sub
